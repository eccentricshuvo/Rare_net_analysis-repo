
module c3540 ( N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, 
        N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, 
        N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, 
        N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, 
        N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, 
        N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, 
        N5231, N5360, N5361 );
  input N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116,
         N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190,
         N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264,
         N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330,
         N343, N349, N350;
  output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815,
         N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231,
         N5360, N5361;
  wire   N26, N323, N538, N5050, N5080, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931;
  assign N1713 = N26;
  assign N3833 = N323;
  assign N5361 = N538;
  assign N5102 = N5050;
  assign N5120 = N5080;

  i1s1 U482 ( .DIN(N179), .Q(n771) );
  hi1s1 U483 ( .DIN(n467), .Q(N538) );
  mxi21s1 U484 ( .DIN1(n467), .DIN2(n468), .SIN(n469), .Q(N5360) );
  and2s1 U485 ( .DIN1(n470), .DIN2(N213), .Q(n469) );
  xor2s1 U486 ( .DIN1(N350), .DIN2(n471), .Q(n468) );
  xor2s1 U487 ( .DIN1(n472), .DIN2(n473), .Q(n467) );
  xnr2s1 U488 ( .DIN1(N5050), .DIN2(n471), .Q(n473) );
  xnr2s1 U489 ( .DIN1(n474), .DIN2(n475), .Q(n471) );
  xor2s1 U490 ( .DIN1(N4815), .DIN2(n476), .Q(n475) );
  xnr2s1 U491 ( .DIN1(N5045), .DIN2(N5121), .Q(n476) );
  xor2s1 U492 ( .DIN1(N5047), .DIN2(n477), .Q(n474) );
  xor2s1 U493 ( .DIN1(N5078), .DIN2(N4944), .Q(n477) );
  nnd3s1 U494 ( .DIN1(n478), .DIN2(N5192), .DIN3(N213), .Q(N5231) );
  oai1112s1 U495 ( .DIN4(n479), .DIN5(n480), .DIN1(n481), .DIN2(n470), .DIN3(
        n472), .Q(n478) );
  hi1s1 U496 ( .DIN(N5080), .Q(n472) );
  hi1s1 U497 ( .DIN(N343), .Q(n470) );
  mxi21s1 U498 ( .DIN1(n482), .DIN2(n483), .SIN(n484), .Q(n480) );
  nnd2s1 U499 ( .DIN1(n485), .DIN2(n486), .Q(n482) );
  or5s1 U500 ( .DIN1(N5078), .DIN2(N5047), .DIN3(N5045), .DIN4(n487), .DIN5(
        n488), .Q(N5192) );
  or5s1 U501 ( .DIN1(N5080), .DIN2(N4815), .DIN3(N5121), .DIN4(n489), .DIN5(
        n490), .Q(n488) );
  hi1s1 U502 ( .DIN(n491), .Q(n490) );
  hi1s1 U503 ( .DIN(n492), .Q(n489) );
  oai13s1 U504 ( .DIN2(n493), .DIN3(n494), .DIN4(n495), .DIN1(n481), .Q(n487)
         );
  oai211s1 U505 ( .DIN1(n496), .DIN2(n497), .DIN3(n479), .DIN4(n498), .Q(n481)
         );
  aoi22s1 U506 ( .DIN1(n499), .DIN2(n500), .DIN3(n501), .DIN4(n502), .Q(n498)
         );
  mxi21s1 U507 ( .DIN1(n503), .DIN2(n504), .SIN(N33), .Q(n499) );
  dsmxc31s1 U508 ( .DIN1(n505), .DIN2(n506), .CLK(n493), .Q(N5121) );
  mxi21s1 U509 ( .DIN1(n507), .DIN2(n508), .SIN(n509), .Q(n506) );
  nnd2s1 U510 ( .DIN1(n510), .DIN2(n511), .Q(n508) );
  oai222s1 U511 ( .DIN1(n512), .DIN2(n495), .DIN3(n513), .DIN4(n514), .DIN5(
        n496), .DIN6(n515), .Q(n505) );
  mxi21s1 U512 ( .DIN1(n516), .DIN2(n517), .SIN(N33), .Q(n512) );
  nnd4s1 U513 ( .DIN1(n518), .DIN2(n519), .DIN3(n520), .DIN4(n521), .Q(n517)
         );
  aoi221s1 U514 ( .DIN1(N107), .DIN2(n522), .DIN3(N97), .DIN4(n523), .DIN5(
        n524), .Q(n521) );
  oai22s1 U515 ( .DIN1(n525), .DIN2(n526), .DIN3(n527), .DIN4(n528), .Q(n524)
         );
  hi1s1 U516 ( .DIN(N303), .Q(n528) );
  aoi22s1 U517 ( .DIN1(N283), .DIN2(n529), .DIN3(N294), .DIN4(n530), .Q(n520)
         );
  nnd4s1 U518 ( .DIN1(n531), .DIN2(n532), .DIN3(n533), .DIN4(n534), .Q(n516)
         );
  aoi22s1 U519 ( .DIN1(N137), .DIN2(n529), .DIN3(N50), .DIN4(n535), .Q(n534)
         );
  aoi22s1 U520 ( .DIN1(N132), .DIN2(n530), .DIN3(N150), .DIN4(n522), .Q(n533)
         );
  aoi22s1 U521 ( .DIN1(N58), .DIN2(n536), .DIN3(N159), .DIN4(n523), .Q(n532)
         );
  aoi22s1 U522 ( .DIN1(N128), .DIN2(n537), .DIN3(N143), .DIN4(n538), .Q(n531)
         );
  mxi21s1 U523 ( .DIN1(n539), .DIN2(n540), .SIN(n479), .Q(N5080) );
  oai322s1 U524 ( .DIN1(n541), .DIN2(N41), .DIN3(n495), .DIN4(N50), .DIN5(n542), .DIN6(n543), .DIN7(n496), .Q(n540) );
  aoi21s1 U525 ( .DIN1(N41), .DIN2(n500), .DIN3(n501), .Q(n542) );
  mxi21s1 U526 ( .DIN1(n544), .DIN2(n545), .SIN(N33), .Q(n541) );
  nnd4s1 U527 ( .DIN1(n546), .DIN2(n547), .DIN3(n548), .DIN4(n549), .Q(n545)
         );
  aoi22s1 U528 ( .DIN1(n529), .DIN2(n550), .DIN3(n535), .DIN4(n513), .Q(n549)
         );
  aoi22s1 U529 ( .DIN1(n530), .DIN2(n526), .DIN3(n522), .DIN4(n551), .Q(n548)
         );
  aoi22s1 U530 ( .DIN1(n536), .DIN2(n502), .DIN3(n523), .DIN4(n552), .Q(n547)
         );
  aoi22s1 U531 ( .DIN1(n537), .DIN2(n553), .DIN3(n538), .DIN4(n554), .Q(n546)
         );
  or3s1 U532 ( .DIN1(n555), .DIN2(n556), .DIN3(n557), .Q(n544) );
  oai221s1 U533 ( .DIN1(n558), .DIN2(N159), .DIN3(n559), .DIN4(N143), .DIN5(
        n560), .Q(n557) );
  hi1s1 U534 ( .DIN(n561), .Q(n560) );
  oai22s1 U535 ( .DIN1(N132), .DIN2(n525), .DIN3(N124), .DIN4(n527), .Q(n561)
         );
  oai22s1 U536 ( .DIN1(n562), .DIN2(N128), .DIN3(n563), .DIN4(N150), .Q(n556)
         );
  oai22s1 U537 ( .DIN1(n564), .DIN2(N125), .DIN3(n565), .DIN4(N137), .Q(n555)
         );
  nnd2s1 U538 ( .DIN1(n566), .DIN2(n567), .Q(n539) );
  oai21s1 U539 ( .DIN1(n509), .DIN2(n484), .DIN3(n507), .Q(n567) );
  and2s1 U540 ( .DIN1(n511), .DIN2(n568), .Q(n507) );
  hi1s1 U541 ( .DIN(n569), .Q(n511) );
  xnr2s1 U542 ( .DIN1(n543), .DIN2(n570), .Q(n566) );
  and2s1 U543 ( .DIN1(n571), .DIN2(n572), .Q(n570) );
  xor2s1 U544 ( .DIN1(n573), .DIN2(n574), .Q(n543) );
  and2s1 U545 ( .DIN1(n575), .DIN2(n576), .Q(n574) );
  oai221s1 U546 ( .DIN1(n577), .DIN2(n578), .DIN3(n579), .DIN4(n580), .DIN5(
        n581), .Q(N5078) );
  aoai1112s1 U547 ( .DIN4(n582), .DIN5(n496), .DIN3(n583), .DIN1(n584), .DIN2(
        n479), .Q(n581) );
  nnd2s1 U548 ( .DIN1(n585), .DIN2(n500), .Q(n584) );
  mxi21s1 U549 ( .DIN1(n586), .DIN2(n587), .SIN(N33), .Q(n585) );
  nnd4s1 U550 ( .DIN1(n588), .DIN2(n589), .DIN3(n590), .DIN4(n591), .Q(n587)
         );
  aoi22s1 U551 ( .DIN1(N311), .DIN2(n529), .DIN3(N116), .DIN4(n535), .Q(n591)
         );
  aoi22s1 U552 ( .DIN1(N317), .DIN2(n530), .DIN3(N294), .DIN4(n522), .Q(n590)
         );
  aoi22s1 U553 ( .DIN1(N107), .DIN2(n536), .DIN3(N283), .DIN4(n523), .Q(n589)
         );
  aoi22s1 U554 ( .DIN1(N322), .DIN2(n537), .DIN3(N303), .DIN4(n538), .Q(n588)
         );
  nnd4s1 U555 ( .DIN1(n592), .DIN2(n593), .DIN3(n594), .DIN4(n595), .Q(n586)
         );
  aoi22s1 U556 ( .DIN1(N159), .DIN2(n529), .DIN3(N77), .DIN4(n535), .Q(n595)
         );
  aoi22s1 U557 ( .DIN1(N150), .DIN2(n530), .DIN3(N58), .DIN4(n522), .Q(n594)
         );
  aoi22s1 U558 ( .DIN1(N87), .DIN2(n536), .DIN3(N68), .DIN4(n523), .Q(n593) );
  aoi22s1 U559 ( .DIN1(N143), .DIN2(n537), .DIN3(N50), .DIN4(n538), .Q(n592)
         );
  aoi21s1 U560 ( .DIN1(n596), .DIN2(n597), .DIN3(n598), .Q(n583) );
  xor2s1 U561 ( .DIN1(n554), .DIN2(n599), .Q(n582) );
  nnd2s1 U562 ( .DIN1(n600), .DIN2(n601), .Q(n599) );
  mxi21s1 U563 ( .DIN1(n602), .DIN2(n603), .SIN(n604), .Q(n578) );
  nor2s1 U564 ( .DIN1(n603), .DIN2(n605), .Q(n602) );
  hi1s1 U565 ( .DIN(n580), .Q(n603) );
  oai21s1 U566 ( .DIN1(n606), .DIN2(n493), .DIN3(n492), .Q(N5050) );
  mxi21s1 U567 ( .DIN1(n607), .DIN2(n483), .SIN(n484), .Q(n492) );
  nnd2s1 U568 ( .DIN1(n608), .DIN2(n571), .Q(n484) );
  mxi21s1 U569 ( .DIN1(n609), .DIN2(n610), .SIN(n497), .Q(n608) );
  aoi21s1 U570 ( .DIN1(n611), .DIN2(n612), .DIN3(n610), .Q(n609) );
  and2s1 U571 ( .DIN1(n485), .DIN2(n510), .Q(n483) );
  oai21s1 U572 ( .DIN1(n485), .DIN2(n577), .DIN3(n568), .Q(n607) );
  nor2s1 U573 ( .DIN1(n509), .DIN2(n569), .Q(n485) );
  oai21s1 U574 ( .DIN1(n613), .DIN2(n614), .DIN3(n615), .Q(n569) );
  xor2s1 U575 ( .DIN1(n616), .DIN2(n515), .Q(n509) );
  oai21s1 U576 ( .DIN1(n613), .DIN2(n617), .DIN3(n618), .Q(n616) );
  aoi222s1 U577 ( .DIN1(n619), .DIN2(n497), .DIN3(n501), .DIN4(N58), .DIN5(
        n500), .DIN6(n620), .Q(n606) );
  dsmxc31s1 U578 ( .DIN1(n504), .DIN2(n503), .CLK(n621), .Q(n620) );
  nnd4s1 U579 ( .DIN1(n622), .DIN2(n623), .DIN3(n624), .DIN4(n625), .Q(n503)
         );
  aoi22s1 U580 ( .DIN1(N132), .DIN2(n529), .DIN3(N159), .DIN4(n535), .Q(n625)
         );
  aoi22s1 U581 ( .DIN1(N128), .DIN2(n530), .DIN3(N143), .DIN4(n522), .Q(n624)
         );
  aoi22s1 U582 ( .DIN1(N50), .DIN2(n536), .DIN3(N150), .DIN4(n523), .Q(n623)
         );
  aoi22s1 U583 ( .DIN1(N125), .DIN2(n537), .DIN3(N137), .DIN4(n538), .Q(n622)
         );
  nnd4s1 U584 ( .DIN1(n626), .DIN2(n627), .DIN3(n628), .DIN4(n629), .Q(n504)
         );
  aoi22s1 U585 ( .DIN1(N116), .DIN2(n529), .DIN3(N77), .DIN4(n535), .Q(n629)
         );
  aoi22s1 U586 ( .DIN1(N283), .DIN2(n530), .DIN3(N97), .DIN4(n522), .Q(n628)
         );
  aoi22s1 U587 ( .DIN1(N68), .DIN2(n536), .DIN3(N87), .DIN4(n523), .Q(n627) );
  aoi22s1 U588 ( .DIN1(N294), .DIN2(n537), .DIN3(N107), .DIN4(n538), .Q(n626)
         );
  hi1s1 U589 ( .DIN(n514), .Q(n501) );
  nnd2s1 U590 ( .DIN1(n495), .DIN2(n496), .Q(n514) );
  nnd2s1 U591 ( .DIN1(n630), .DIN2(n631), .Q(N5047) );
  oai211s1 U592 ( .DIN1(n632), .DIN2(n633), .DIN3(n479), .DIN4(n634), .Q(n631)
         );
  aoi22s1 U593 ( .DIN1(n635), .DIN2(n500), .DIN3(n598), .DIN4(n636), .Q(n634)
         );
  oai21s1 U594 ( .DIN1(n637), .DIN2(n638), .DIN3(n639), .Q(n636) );
  mxi21s1 U595 ( .DIN1(n640), .DIN2(n641), .SIN(n642), .Q(n639) );
  nor2s1 U596 ( .DIN1(N107), .DIN2(n601), .Q(n641) );
  mxi21s1 U597 ( .DIN1(n643), .DIN2(n644), .SIN(N45), .Q(n637) );
  oai1112s1 U598 ( .DIN4(n513), .DIN5(n552), .DIN1(n645), .DIN2(N58), .DIN3(
        n646), .Q(n643) );
  hi1s1 U599 ( .DIN(n640), .Q(n645) );
  mxi21s1 U600 ( .DIN1(n647), .DIN2(n648), .SIN(N33), .Q(n635) );
  nnd4s1 U601 ( .DIN1(n649), .DIN2(n650), .DIN3(n651), .DIN4(n652), .Q(n648)
         );
  aoi22s1 U602 ( .DIN1(N317), .DIN2(n529), .DIN3(N283), .DIN4(n535), .Q(n652)
         );
  aoi22s1 U603 ( .DIN1(N322), .DIN2(n530), .DIN3(N303), .DIN4(n522), .Q(n651)
         );
  aoi22s1 U604 ( .DIN1(N326), .DIN2(n537), .DIN3(N294), .DIN4(n523), .Q(n650)
         );
  aoi22s1 U605 ( .DIN1(N116), .DIN2(n536), .DIN3(N311), .DIN4(n538), .Q(n649)
         );
  oai1112s1 U606 ( .DIN4(n558), .DIN5(n554), .DIN1(n519), .DIN2(n653), .DIN3(
        n654), .Q(n647) );
  aoi221s1 U607 ( .DIN1(N58), .DIN2(n538), .DIN3(N50), .DIN4(n529), .DIN5(n655), .Q(n654) );
  oai22s1 U608 ( .DIN1(n564), .DIN2(n656), .DIN3(n565), .DIN4(n513), .Q(n655)
         );
  aoi22s1 U609 ( .DIN1(N77), .DIN2(n523), .DIN3(N150), .DIN4(n537), .Q(n653)
         );
  nnd2s1 U610 ( .DIN1(N87), .DIN2(n535), .Q(n519) );
  mxi21s1 U611 ( .DIN1(n657), .DIN2(n658), .SIN(n604), .Q(n630) );
  nor2s1 U612 ( .DIN1(n577), .DIN2(n605), .Q(n658) );
  oai21s1 U613 ( .DIN1(n659), .DIN2(n660), .DIN3(n661), .Q(N5045) );
  aoai1112s1 U614 ( .DIN4(n662), .DIN5(n642), .DIN3(n663), .DIN1(n479), .DIN2(
        n664), .Q(n661) );
  aoi22s1 U615 ( .DIN1(n665), .DIN2(n500), .DIN3(n666), .DIN4(n597), .Q(n664)
         );
  mxi21s1 U616 ( .DIN1(n667), .DIN2(n668), .SIN(N33), .Q(n665) );
  nnd4s1 U617 ( .DIN1(n669), .DIN2(n670), .DIN3(n671), .DIN4(n672), .Q(n668)
         );
  aoi22s1 U618 ( .DIN1(N97), .DIN2(n536), .DIN3(N116), .DIN4(n523), .Q(n672)
         );
  aoi22s1 U619 ( .DIN1(N317), .DIN2(n537), .DIN3(N294), .DIN4(n538), .Q(n671)
         );
  aoi22s1 U620 ( .DIN1(N303), .DIN2(n529), .DIN3(N311), .DIN4(n530), .Q(n670)
         );
  aoi22s1 U621 ( .DIN1(N283), .DIN2(n522), .DIN3(N107), .DIN4(n535), .Q(n669)
         );
  oai1112s1 U622 ( .DIN4(n562), .DIN5(n673), .DIN1(n518), .DIN2(n674), .DIN3(
        n675), .Q(n667) );
  aoi221s1 U623 ( .DIN1(N58), .DIN2(n523), .DIN3(N159), .DIN4(n538), .DIN5(
        n676), .Q(n675) );
  oai22s1 U624 ( .DIN1(n527), .DIN2(n677), .DIN3(n565), .DIN4(n646), .Q(n676)
         );
  hi1s1 U625 ( .DIN(N137), .Q(n677) );
  aoi22s1 U626 ( .DIN1(N68), .DIN2(n535), .DIN3(N143), .DIN4(n530), .Q(n674)
         );
  nnd2s1 U627 ( .DIN1(N77), .DIN2(n536), .Q(n518) );
  mxi21s1 U628 ( .DIN1(n551), .DIN2(n678), .SIN(n601), .Q(n662) );
  oai13s1 U629 ( .DIN2(n666), .DIN3(n679), .DIN4(n680), .DIN1(n681), .Q(n660)
         );
  oai13s1 U630 ( .DIN2(n580), .DIN3(n604), .DIN4(n577), .DIN1(n579), .Q(n681)
         );
  hi1s1 U631 ( .DIN(n657), .Q(n579) );
  oai21s1 U632 ( .DIN1(n613), .DIN2(n577), .DIN3(n568), .Q(n657) );
  aoi13s1 U633 ( .DIN2(N13), .DIN3(n682), .DIN4(N45), .DIN1(n683), .Q(n568) );
  xor2s1 U634 ( .DIN1(n684), .DIN2(n685), .Q(n604) );
  nor2s1 U635 ( .DIN1(n679), .DIN2(n686), .Q(n685) );
  nnd2s1 U636 ( .DIN1(n687), .DIN2(n688), .Q(n684) );
  hi1s1 U637 ( .DIN(n689), .Q(n688) );
  aoi21s1 U638 ( .DIN1(n690), .DIN2(N330), .DIN3(n632), .Q(n689) );
  xor2s1 U639 ( .DIN1(n596), .DIN2(N4589), .Q(n580) );
  mxi21s1 U640 ( .DIN1(n691), .DIN2(n692), .SIN(n693), .Q(n659) );
  nor2s1 U641 ( .DIN1(n596), .DIN2(n687), .Q(n693) );
  xor2s1 U642 ( .DIN1(n694), .DIN2(n666), .Q(n692) );
  aoi22s1 U643 ( .DIN1(n695), .DIN2(n666), .DIN3(n694), .DIN4(n696), .Q(n691)
         );
  nor2s1 U644 ( .DIN1(n697), .DIN2(n698), .Q(n694) );
  dsmxc31s1 U645 ( .DIN1(n698), .DIN2(n680), .CLK(n697), .Q(n695) );
  hi1s1 U646 ( .DIN(n699), .Q(n680) );
  oai21s1 U647 ( .DIN1(n700), .DIN2(n596), .DIN3(n701), .Q(n699) );
  xor2s1 U648 ( .DIN1(n702), .DIN2(n703), .Q(n596) );
  nnd2s1 U649 ( .DIN1(n679), .DIN2(n704), .Q(n702) );
  oai13s1 U650 ( .DIN2(n705), .DIN3(n706), .DIN4(n526), .DIN1(n707), .Q(N5002)
         );
  mxi21s1 U651 ( .DIN1(n708), .DIN2(n709), .SIN(n710), .Q(n707) );
  nor2s1 U652 ( .DIN1(n711), .DIN2(n712), .Q(n709) );
  xor2s1 U653 ( .DIN1(n713), .DIN2(n714), .Q(n712) );
  xnr2s1 U654 ( .DIN1(n572), .DIN2(n715), .Q(n714) );
  oai21s1 U655 ( .DIN1(n614), .DIN2(n716), .DIN3(n615), .Q(n715) );
  aoi22s1 U656 ( .DIN1(n610), .DIN2(n497), .DIN3(n717), .DIN4(n718), .Q(n572)
         );
  hi1s1 U657 ( .DIN(n719), .Q(n718) );
  oai222s1 U658 ( .DIN1(n515), .DIN2(n618), .DIN3(n720), .DIN4(n716), .DIN5(
        n679), .DIN6(n721), .Q(n610) );
  hi1s1 U659 ( .DIN(n611), .Q(n720) );
  mxi21s1 U660 ( .DIN1(n722), .DIN2(n723), .SIN(n614), .Q(n713) );
  hi1s1 U661 ( .DIN(n571), .Q(n723) );
  nnd3s1 U662 ( .DIN1(n612), .DIN2(n497), .DIN3(n611), .Q(n571) );
  hi1s1 U663 ( .DIN(n724), .Q(n612) );
  aoi21s1 U664 ( .DIN1(n611), .DIN2(n497), .DIN3(n724), .Q(n722) );
  xor2s1 U665 ( .DIN1(n725), .DIN2(n726), .Q(n497) );
  nnd2s1 U666 ( .DIN1(n576), .DIN2(n727), .Q(n725) );
  nor2s1 U667 ( .DIN1(n617), .DIN2(n515), .Q(n611) );
  nnd2s1 U668 ( .DIN1(n728), .DIN2(n729), .Q(n515) );
  mxi21s1 U669 ( .DIN1(n730), .DIN2(n731), .SIN(n679), .Q(n728) );
  nor2s1 U670 ( .DIN1(n732), .DIN2(n733), .Q(n731) );
  hi1s1 U671 ( .DIN(n705), .Q(n711) );
  oai22s1 U672 ( .DIN1(N50), .DIN2(n513), .DIN3(n552), .DIN4(n734), .Q(n708)
         );
  mxi21s1 U673 ( .DIN1(N68), .DIN2(n735), .SIN(N58), .Q(n734) );
  nor2s1 U674 ( .DIN1(N68), .DIN2(n646), .Q(n735) );
  oai13s1 U675 ( .DIN2(n493), .DIN3(n494), .DIN4(n495), .DIN1(n491), .Q(N4944)
         );
  mxi21s1 U676 ( .DIN1(n736), .DIN2(n737), .SIN(n479), .Q(n491) );
  hi1s1 U677 ( .DIN(n493), .Q(n479) );
  nor2s1 U678 ( .DIN1(n500), .DIN2(n738), .Q(n737) );
  dsmxc31s1 U679 ( .DIN1(n617), .DIN2(n552), .CLK(n496), .Q(n738) );
  xor2s1 U680 ( .DIN1(n617), .DIN2(n613), .Q(n736) );
  hi1s1 U681 ( .DIN(n605), .Q(n613) );
  nnd2s1 U682 ( .DIN1(n739), .DIN2(n618), .Q(n617) );
  nnd2s1 U683 ( .DIN1(n740), .DIN2(n697), .Q(n618) );
  mxi21s1 U684 ( .DIN1(n741), .DIN2(n742), .SIN(n743), .Q(n739) );
  nor2s1 U685 ( .DIN1(n740), .DIN2(n697), .Q(n741) );
  mxi21s1 U686 ( .DIN1(n744), .DIN2(n745), .SIN(N33), .Q(n494) );
  nnd4s1 U687 ( .DIN1(n746), .DIN2(n747), .DIN3(n748), .DIN4(n749), .Q(n745)
         );
  aoi22s1 U688 ( .DIN1(N294), .DIN2(n529), .DIN3(N97), .DIN4(n535), .Q(n749)
         );
  aoi22s1 U689 ( .DIN1(N303), .DIN2(n530), .DIN3(N116), .DIN4(n522), .Q(n748)
         );
  aoi22s1 U690 ( .DIN1(N87), .DIN2(n536), .DIN3(N107), .DIN4(n523), .Q(n747)
         );
  aoi22s1 U691 ( .DIN1(N311), .DIN2(n537), .DIN3(N283), .DIN4(n538), .Q(n746)
         );
  nnd4s1 U692 ( .DIN1(n750), .DIN2(n751), .DIN3(n752), .DIN4(n753), .Q(n744)
         );
  aoi22s1 U693 ( .DIN1(N143), .DIN2(n529), .DIN3(N58), .DIN4(n535), .Q(n753)
         );
  aoi22s1 U694 ( .DIN1(N137), .DIN2(n530), .DIN3(N159), .DIN4(n522), .Q(n752)
         );
  aoi22s1 U695 ( .DIN1(N68), .DIN2(n536), .DIN3(N50), .DIN4(n523), .Q(n751) );
  aoi22s1 U696 ( .DIN1(N132), .DIN2(n537), .DIN3(N150), .DIN4(n538), .Q(n750)
         );
  dsmxc31s1 U697 ( .DIN1(n754), .DIN2(n755), .CLK(n493), .Q(N4815) );
  nnd2s1 U698 ( .DIN1(n486), .DIN2(n577), .Q(n493) );
  nnd2s1 U699 ( .DIN1(n710), .DIN2(n756), .Q(n486) );
  oai21s1 U700 ( .DIN1(N20), .DIN2(n757), .DIN3(N1), .Q(n756) );
  xor2s1 U701 ( .DIN1(N330), .DIN2(n690), .Q(n755) );
  aoi222s1 U702 ( .DIN1(n598), .DIN2(n758), .DIN3(n759), .DIN4(n500), .DIN5(
        n760), .DIN6(n597), .Q(n754) );
  hi1s1 U703 ( .DIN(n633), .Q(n597) );
  hi1s1 U704 ( .DIN(n690), .Q(n760) );
  hi1s1 U705 ( .DIN(n495), .Q(n500) );
  mxi21s1 U706 ( .DIN1(n761), .DIN2(n762), .SIN(N33), .Q(n759) );
  nnd4s1 U707 ( .DIN1(n763), .DIN2(n764), .DIN3(n765), .DIN4(n766), .Q(n762)
         );
  aoi22s1 U708 ( .DIN1(N283), .DIN2(n536), .DIN3(N303), .DIN4(n523), .Q(n766)
         );
  aoi22s1 U709 ( .DIN1(N329), .DIN2(n537), .DIN3(N317), .DIN4(n538), .Q(n765)
         );
  aoi22s1 U710 ( .DIN1(N322), .DIN2(n529), .DIN3(N311), .DIN4(n522), .Q(n764)
         );
  aoi22s1 U711 ( .DIN1(N326), .DIN2(n530), .DIN3(N294), .DIN4(n535), .Q(n763)
         );
  nnd4s1 U712 ( .DIN1(n767), .DIN2(n768), .DIN3(n769), .DIN4(n770), .Q(n761)
         );
  aoi22s1 U713 ( .DIN1(N107), .DIN2(n536), .DIN3(N87), .DIN4(n523), .Q(n770)
         );
  hi1s1 U714 ( .DIN(n559), .Q(n523) );
  nnd3s1 U715 ( .DIN1(N190), .DIN2(n771), .DIN3(n772), .Q(n559) );
  hi1s1 U716 ( .DIN(n558), .Q(n536) );
  nnd3s1 U717 ( .DIN1(n771), .DIN2(n773), .DIN3(n772), .Q(n558) );
  aoi22s1 U718 ( .DIN1(N159), .DIN2(n537), .DIN3(N68), .DIN4(n538), .Q(n769)
         );
  hi1s1 U719 ( .DIN(n525), .Q(n538) );
  nnd3s1 U720 ( .DIN1(N179), .DIN2(n773), .DIN3(n772), .Q(n525) );
  hi1s1 U721 ( .DIN(n527), .Q(n537) );
  nnd2s1 U722 ( .DIN1(n774), .DIN2(n771), .Q(n527) );
  aoi22s1 U723 ( .DIN1(N50), .DIN2(n530), .DIN3(N77), .DIN4(n522), .Q(n768) );
  hi1s1 U724 ( .DIN(n565), .Q(n522) );
  nnd2s1 U725 ( .DIN1(n774), .DIN2(N179), .Q(n565) );
  and3s1 U726 ( .DIN1(n773), .DIN2(n775), .DIN3(N20), .Q(n774) );
  hi1s1 U727 ( .DIN(n564), .Q(n530) );
  nnd3s1 U728 ( .DIN1(N179), .DIN2(N190), .DIN3(n772), .Q(n564) );
  nor2s1 U729 ( .DIN1(n775), .DIN2(n682), .Q(n772) );
  aoi22s1 U730 ( .DIN1(N58), .DIN2(n529), .DIN3(N97), .DIN4(n535), .Q(n767) );
  hi1s1 U731 ( .DIN(n563), .Q(n535) );
  aoi21s1 U732 ( .DIN1(n771), .DIN2(n776), .DIN3(n682), .Q(n563) );
  hi1s1 U733 ( .DIN(n562), .Q(n529) );
  nnd3s1 U734 ( .DIN1(n776), .DIN2(N20), .DIN3(N179), .Q(n562) );
  nor2s1 U735 ( .DIN1(n773), .DIN2(N200), .Q(n776) );
  oai21s1 U736 ( .DIN1(n777), .DIN2(n638), .DIN3(n778), .Q(n758) );
  mxi21s1 U737 ( .DIN1(N1947), .DIN2(n779), .SIN(n642), .Q(n778) );
  nnd2s1 U738 ( .DIN1(n780), .DIN2(n621), .Q(n642) );
  nor2s1 U739 ( .DIN1(N116), .DIN2(n601), .Q(n779) );
  hi1s1 U740 ( .DIN(n638), .Q(n601) );
  nnd2s1 U741 ( .DIN1(N33), .DIN2(n780), .Q(n638) );
  mxi21s1 U742 ( .DIN1(n781), .DIN2(n782), .SIN(N45), .Q(n777) );
  hi1s1 U743 ( .DIN(n663), .Q(n598) );
  nnd2s1 U744 ( .DIN1(n633), .DIN2(n495), .Q(n663) );
  oai21s1 U745 ( .DIN1(N169), .DIN2(n682), .DIN3(n783), .Q(n495) );
  nnd2s1 U746 ( .DIN1(n619), .DIN2(n682), .Q(n633) );
  oai21s1 U747 ( .DIN1(n577), .DIN2(n781), .DIN3(n784), .Q(N4667) );
  mxi21s1 U748 ( .DIN1(n605), .DIN2(n785), .SIN(N1), .Q(n784) );
  nor2s1 U749 ( .DIN1(n510), .DIN2(n640), .Q(n785) );
  nnd3s1 U750 ( .DIN1(n526), .DIN2(n554), .DIN3(n786), .Q(n640) );
  hi1s1 U751 ( .DIN(n577), .Q(n510) );
  nnd2s1 U752 ( .DIN1(n716), .DIN2(n724), .Q(n605) );
  nnd2s1 U753 ( .DIN1(n787), .DIN2(N330), .Q(n724) );
  mxi21s1 U754 ( .DIN1(n788), .DIN2(n789), .SIN(n679), .Q(n787) );
  oai211s1 U755 ( .DIN1(N179), .DIN2(n790), .DIN3(n791), .DIN4(n792), .Q(n789)
         );
  mxi21s1 U756 ( .DIN1(n790), .DIN2(n793), .SIN(n794), .Q(n792) );
  mxi21s1 U757 ( .DIN1(N179), .DIN2(n795), .SIN(n796), .Q(n791) );
  nnd4s1 U758 ( .DIN1(n703), .DIN2(n797), .DIN3(n798), .DIN4(n696), .Q(n788)
         );
  hi1s1 U759 ( .DIN(n666), .Q(n696) );
  aoi21s1 U760 ( .DIN1(n799), .DIN2(n800), .DIN3(n801), .Q(n798) );
  nnd2s1 U761 ( .DIN1(n802), .DIN2(n697), .Q(n716) );
  nnd2s1 U762 ( .DIN1(n780), .DIN2(n803), .Q(n577) );
  oai21s1 U763 ( .DIN1(n679), .DIN2(n700), .DIN3(n687), .Q(N4589) );
  nnd3s1 U764 ( .DIN1(n632), .DIN2(n690), .DIN3(N330), .Q(n687) );
  oai21s1 U765 ( .DIN1(n800), .DIN2(n804), .DIN3(n805), .Q(n690) );
  mxi21s1 U766 ( .DIN1(n806), .DIN2(n801), .SIN(n679), .Q(n805) );
  nor2s1 U767 ( .DIN1(n799), .DIN2(n807), .Q(n806) );
  hi1s1 U768 ( .DIN(n804), .Q(n799) );
  aoi21s1 U769 ( .DIN1(n632), .DIN2(n801), .DIN3(n808), .Q(n700) );
  hi1s1 U770 ( .DIN(n809), .Q(n808) );
  hi1s1 U771 ( .DIN(n686), .Q(n801) );
  xnr2s1 U772 ( .DIN1(n810), .DIN2(n797), .Q(n632) );
  hi1s1 U773 ( .DIN(n811), .Q(n797) );
  nnd2s1 U774 ( .DIN1(n679), .DIN2(n812), .Q(n810) );
  hi1s1 U775 ( .DIN(n697), .Q(n679) );
  nnd2s1 U776 ( .DIN1(N343), .DIN2(n576), .Q(n697) );
  hi1s1 U777 ( .DIN(n717), .Q(n576) );
  nnd4s1 U778 ( .DIN1(N213), .DIN2(N13), .DIN3(n683), .DIN4(n682), .Q(n717) );
  oai21s1 U779 ( .DIN1(n813), .DIN2(n614), .DIN3(n615), .Q(N4145) );
  aoi22s1 U780 ( .DIN1(n814), .DIN2(n573), .DIN3(n575), .DIN4(n815), .Q(n615)
         );
  mxi21s1 U781 ( .DIN1(n771), .DIN2(n816), .SIN(n817), .Q(n815) );
  oai211s1 U782 ( .DIN1(n818), .DIN2(n673), .DIN3(n819), .DIN4(n820), .Q(n575)
         );
  aoi22s1 U783 ( .DIN1(N58), .DIN2(n821), .DIN3(N68), .DIN4(n822), .Q(n820) );
  hi1s1 U784 ( .DIN(n823), .Q(n821) );
  mxi21s1 U785 ( .DIN1(n824), .DIN2(n825), .SIN(N50), .Q(n819) );
  hi1s1 U786 ( .DIN(N150), .Q(n673) );
  oai21s1 U787 ( .DIN1(n726), .DIN2(n826), .DIN3(n719), .Q(n814) );
  aoi21s1 U788 ( .DIN1(n729), .DIN2(n740), .DIN3(n730), .Q(n826) );
  hi1s1 U789 ( .DIN(n721), .Q(n730) );
  hi1s1 U790 ( .DIN(n827), .Q(n740) );
  hi1s1 U791 ( .DIN(n802), .Q(n813) );
  oai22s1 U792 ( .DIN1(n698), .DIN2(n828), .DIN3(n829), .DIN4(n666), .Q(n802)
         );
  aoi21s1 U793 ( .DIN1(n703), .DIN2(n830), .DIN3(n831), .Q(n829) );
  hi1s1 U794 ( .DIN(n701), .Q(n831) );
  oai21s1 U795 ( .DIN1(n811), .DIN2(n686), .DIN3(n809), .Q(n830) );
  nnd2s1 U796 ( .DIN1(n807), .DIN2(n804), .Q(n686) );
  hi1s1 U797 ( .DIN(n832), .Q(n703) );
  mxi21s1 U798 ( .DIN1(N169), .DIN2(N179), .SIN(n796), .Q(n828) );
  aoi211s1 U799 ( .DIN1(N68), .DIN2(n833), .DIN3(n834), .DIN4(n835), .Q(n698)
         );
  mxi21s1 U800 ( .DIN1(n836), .DIN2(n837), .SIN(n551), .Q(n834) );
  nor5s1 U801 ( .DIN1(n614), .DIN2(n838), .DIN3(n832), .DIN4(n666), .DIN5(n811), .Q(N4028) );
  oai21s1 U802 ( .DIN1(n812), .DIN2(n839), .DIN3(n809), .Q(n811) );
  nnd2s1 U803 ( .DIN1(n840), .DIN2(n812), .Q(n809) );
  mxi21s1 U804 ( .DIN1(n771), .DIN2(n816), .SIN(n794), .Q(n840) );
  mxi21s1 U805 ( .DIN1(n773), .DIN2(n775), .SIN(n794), .Q(n839) );
  oai211s1 U806 ( .DIN1(n841), .DIN2(n842), .DIN3(n843), .DIN4(n844), .Q(n794)
         );
  aoi22s1 U807 ( .DIN1(N264), .DIN2(n845), .DIN3(N294), .DIN4(n846), .Q(n844)
         );
  mxi21s1 U808 ( .DIN1(N250), .DIN2(N257), .SIN(N349), .Q(n842) );
  oai221s1 U809 ( .DIN1(n847), .DIN2(n526), .DIN3(n818), .DIN4(n551), .DIN5(
        n848), .Q(n812) );
  mxi21s1 U810 ( .DIN1(n849), .DIN2(n850), .SIN(N107), .Q(n848) );
  hi1s1 U811 ( .DIN(N116), .Q(n526) );
  mxi41s1 U812 ( .DIN1(n816), .DIN2(n771), .DIN3(N200), .DIN4(N190), .SIN0(
        n796), .SIN1(n851), .Q(n666) );
  aoi211s1 U813 ( .DIN1(n833), .DIN2(N68), .DIN3(n835), .DIN4(n852), .Q(n851)
         );
  mxi21s1 U814 ( .DIN1(n837), .DIN2(n836), .SIN(N87), .Q(n852) );
  oai22s1 U815 ( .DIN1(n853), .DIN2(n786), .DIN3(n554), .DIN4(n823), .Q(n835)
         );
  aoi221s1 U816 ( .DIN1(n854), .DIN2(n855), .DIN3(n846), .DIN4(N116), .DIN5(
        n856), .Q(n796) );
  dsmxc31s1 U817 ( .DIN1(n857), .DIN2(N274), .CLK(n858), .Q(n856) );
  and2s1 U818 ( .DIN1(n859), .DIN2(N250), .Q(n857) );
  dsmxc31s1 U819 ( .DIN1(N238), .DIN2(N244), .CLK(N349), .Q(n855) );
  oai21s1 U820 ( .DIN1(n704), .DIN2(n860), .DIN3(n701), .Q(n832) );
  nnd2s1 U821 ( .DIN1(n861), .DIN2(n704), .Q(n701) );
  mxi21s1 U822 ( .DIN1(n771), .DIN2(n816), .SIN(n790), .Q(n861) );
  mxi21s1 U823 ( .DIN1(n773), .DIN2(n775), .SIN(n790), .Q(n860) );
  oai211s1 U824 ( .DIN1(n841), .DIN2(n862), .DIN3(n843), .DIN4(n863), .Q(n790)
         );
  aoi22s1 U825 ( .DIN1(N257), .DIN2(n845), .DIN3(N283), .DIN4(n846), .Q(n863)
         );
  mxi21s1 U826 ( .DIN1(N244), .DIN2(N250), .SIN(N349), .Q(n862) );
  oai211s1 U827 ( .DIN1(n818), .DIN2(n552), .DIN3(n864), .DIN4(n865), .Q(n704)
         );
  aoi22s1 U828 ( .DIN1(N107), .DIN2(n866), .DIN3(n706), .DIN4(n822), .Q(n865)
         );
  xor2s1 U829 ( .DIN1(n550), .DIN2(N97), .Q(n706) );
  mxi21s1 U830 ( .DIN1(n824), .DIN2(n850), .SIN(N97), .Q(n864) );
  hi1s1 U831 ( .DIN(n836), .Q(n850) );
  dsmxc31s1 U832 ( .DIN1(n800), .DIN2(n807), .CLK(n804), .Q(n838) );
  oai221s1 U833 ( .DIN1(n847), .DIN2(n553), .DIN3(n818), .DIN4(n554), .DIN5(
        n867), .Q(n804) );
  mxi21s1 U834 ( .DIN1(n824), .DIN2(n868), .SIN(N116), .Q(n867) );
  nnd2s1 U835 ( .DIN1(n853), .DIN2(n836), .Q(n868) );
  oai21s1 U836 ( .DIN1(N1), .DIN2(n621), .DIN3(n869), .Q(n836) );
  hi1s1 U837 ( .DIN(N97), .Q(n554) );
  hi1s1 U838 ( .DIN(N283), .Q(n553) );
  mxi21s1 U839 ( .DIN1(n816), .DIN2(n771), .SIN(n793), .Q(n807) );
  mxi21s1 U840 ( .DIN1(N200), .DIN2(N190), .SIN(n793), .Q(n800) );
  hi1s1 U841 ( .DIN(n795), .Q(n793) );
  oai211s1 U842 ( .DIN1(n841), .DIN2(n870), .DIN3(n843), .DIN4(n871), .Q(n795)
         );
  aoi22s1 U843 ( .DIN1(N270), .DIN2(n845), .DIN3(N303), .DIN4(n846), .Q(n871)
         );
  nor2s1 U844 ( .DIN1(n872), .DIN2(n873), .Q(n845) );
  nnd2s1 U845 ( .DIN1(n872), .DIN2(N274), .Q(n843) );
  and2s1 U846 ( .DIN1(n858), .DIN2(n803), .Q(n872) );
  nor2s1 U847 ( .DIN1(n757), .DIN2(N1), .Q(n858) );
  mxi21s1 U848 ( .DIN1(N257), .DIN2(N264), .SIN(N349), .Q(n870) );
  nnd4s1 U849 ( .DIN1(n827), .DIN2(n721), .DIN3(n729), .DIN4(n874), .Q(n614)
         );
  aoi211s1 U850 ( .DIN1(n743), .DIN2(n742), .DIN3(n726), .DIN4(n875), .Q(n874)
         );
  hi1s1 U851 ( .DIN(n573), .Q(n875) );
  mxi41s1 U852 ( .DIN1(N179), .DIN2(N169), .DIN3(n773), .DIN4(n775), .SIN0(
        n817), .SIN1(n876), .Q(n573) );
  aoi211s1 U853 ( .DIN1(N150), .DIN2(n833), .DIN3(n877), .DIN4(n878), .Q(n876)
         );
  mxi21s1 U854 ( .DIN1(n837), .DIN2(n879), .SIN(N50), .Q(n878) );
  oai22s1 U855 ( .DIN1(n853), .DIN2(n513), .DIN3(n823), .DIN4(n502), .Q(n877)
         );
  aoi21s1 U856 ( .DIN1(N33), .DIN2(n880), .DIN3(n822), .Q(n823) );
  hi1s1 U857 ( .DIN(n818), .Q(n833) );
  oai211s1 U858 ( .DIN1(n841), .DIN2(n881), .DIN3(n882), .DIN4(n883), .Q(n817)
         );
  aoi22s1 U859 ( .DIN1(N226), .DIN2(n884), .DIN3(N77), .DIN4(n846), .Q(n883)
         );
  mxi21s1 U860 ( .DIN1(N222), .DIN2(N223), .SIN(N349), .Q(n881) );
  oai21s1 U861 ( .DIN1(n727), .DIN2(n885), .DIN3(n719), .Q(n726) );
  nnd2s1 U862 ( .DIN1(n886), .DIN2(n727), .Q(n719) );
  mxi21s1 U863 ( .DIN1(n771), .DIN2(n816), .SIN(n887), .Q(n886) );
  mxi21s1 U864 ( .DIN1(n773), .DIN2(n775), .SIN(n887), .Q(n885) );
  oai211s1 U865 ( .DIN1(n888), .DIN2(n889), .DIN3(n882), .DIN4(n890), .Q(n887)
         );
  aoi22s1 U866 ( .DIN1(N87), .DIN2(n846), .DIN3(n891), .DIN4(n854), .Q(n890)
         );
  dsmxc31s1 U867 ( .DIN1(N223), .DIN2(N226), .CLK(N349), .Q(n891) );
  hi1s1 U868 ( .DIN(N200), .Q(n775) );
  hi1s1 U869 ( .DIN(N190), .Q(n773) );
  oai211s1 U870 ( .DIN1(n818), .DIN2(n656), .DIN3(n892), .DIN4(n893), .Q(n727)
         );
  aoi22s1 U871 ( .DIN1(n866), .DIN2(N68), .DIN3(n822), .DIN4(n894), .Q(n893)
         );
  hi1s1 U872 ( .DIN(n847), .Q(n866) );
  mxi21s1 U873 ( .DIN1(n824), .DIN2(n895), .SIN(N58), .Q(n892) );
  hi1s1 U874 ( .DIN(N159), .Q(n656) );
  mxi21s1 U875 ( .DIN1(N190), .DIN2(N200), .SIN(n896), .Q(n742) );
  hi1s1 U876 ( .DIN(n897), .Q(n743) );
  nnd2s1 U877 ( .DIN1(n898), .DIN2(n732), .Q(n729) );
  hi1s1 U878 ( .DIN(n899), .Q(n732) );
  mxi21s1 U879 ( .DIN1(N190), .DIN2(N200), .SIN(n900), .Q(n898) );
  nnd2s1 U880 ( .DIN1(n733), .DIN2(n899), .Q(n721) );
  oai221s1 U881 ( .DIN1(n552), .DIN2(n847), .DIN3(n818), .DIN4(n646), .DIN5(
        n901), .Q(n899) );
  mxi21s1 U882 ( .DIN1(n849), .DIN2(n895), .SIN(N68), .Q(n901) );
  nnd2s1 U883 ( .DIN1(n853), .DIN2(n837), .Q(n849) );
  hi1s1 U884 ( .DIN(n824), .Q(n837) );
  hi1s1 U885 ( .DIN(N77), .Q(n552) );
  mxi21s1 U886 ( .DIN1(n771), .DIN2(n816), .SIN(n900), .Q(n733) );
  oai211s1 U887 ( .DIN1(n888), .DIN2(n902), .DIN3(n882), .DIN4(n903), .Q(n900)
         );
  aoi22s1 U888 ( .DIN1(N97), .DIN2(n846), .DIN3(n904), .DIN4(n854), .Q(n903)
         );
  hi1s1 U889 ( .DIN(n841), .Q(n854) );
  dsmxc31s1 U890 ( .DIN1(N226), .DIN2(N232), .CLK(N349), .Q(n904) );
  hi1s1 U891 ( .DIN(n884), .Q(n888) );
  nnd2s1 U892 ( .DIN1(n905), .DIN2(n897), .Q(n827) );
  oai221s1 U893 ( .DIN1(n847), .DIN2(n551), .DIN3(n502), .DIN4(n818), .DIN5(
        n906), .Q(n897) );
  mxi21s1 U894 ( .DIN1(n824), .DIN2(n825), .SIN(N77), .Q(n906) );
  hi1s1 U895 ( .DIN(n879), .Q(n825) );
  nor2s1 U896 ( .DIN1(n822), .DIN2(n895), .Q(n879) );
  and2s1 U897 ( .DIN1(n869), .DIN2(n907), .Q(n895) );
  nor2s1 U898 ( .DIN1(n824), .DIN2(n880), .Q(n869) );
  hi1s1 U899 ( .DIN(n853), .Q(n822) );
  nnd2s1 U900 ( .DIN1(n880), .DIN2(N20), .Q(n853) );
  nor2s1 U901 ( .DIN1(n907), .DIN2(n908), .Q(n824) );
  nnd2s1 U902 ( .DIN1(N20), .DIN2(n683), .Q(n907) );
  nnd3s1 U903 ( .DIN1(n682), .DIN2(n621), .DIN3(n880), .Q(n818) );
  nnd3s1 U904 ( .DIN1(N33), .DIN2(n682), .DIN3(n880), .Q(n847) );
  aoi211s1 U905 ( .DIN1(n908), .DIN2(n682), .DIN3(n619), .DIN4(n683), .Q(n880)
         );
  hi1s1 U906 ( .DIN(n496), .Q(n619) );
  nnd2s1 U907 ( .DIN1(n908), .DIN2(n621), .Q(n496) );
  mxi21s1 U908 ( .DIN1(n771), .DIN2(n816), .SIN(n896), .Q(n905) );
  oai211s1 U909 ( .DIN1(n841), .DIN2(n909), .DIN3(n882), .DIN4(n910), .Q(n896)
         );
  aoi22s1 U910 ( .DIN1(N244), .DIN2(n884), .DIN3(N107), .DIN4(n846), .Q(n910)
         );
  nor2s1 U911 ( .DIN1(n859), .DIN2(n621), .Q(n846) );
  nor2s1 U912 ( .DIN1(n873), .DIN2(n911), .Q(n884) );
  nnd2s1 U913 ( .DIN1(N274), .DIN2(n911), .Q(n882) );
  aoi21s1 U914 ( .DIN1(n757), .DIN2(n803), .DIN3(N1), .Q(n911) );
  hi1s1 U915 ( .DIN(N45), .Q(n757) );
  mxi21s1 U916 ( .DIN1(N232), .DIN2(N238), .SIN(N349), .Q(n909) );
  nnd2s1 U917 ( .DIN1(n873), .DIN2(n621), .Q(n841) );
  hi1s1 U918 ( .DIN(n859), .Q(n873) );
  oai21s1 U919 ( .DIN1(n621), .DIN2(n803), .DIN3(n783), .Q(n859) );
  hi1s1 U920 ( .DIN(N41), .Q(n803) );
  hi1s1 U921 ( .DIN(N33), .Q(n621) );
  hi1s1 U922 ( .DIN(N169), .Q(n816) );
  xor2s1 U923 ( .DIN1(n782), .DIN2(n912), .Q(N3987) );
  xor2s1 U924 ( .DIN1(N97), .DIN2(n600), .Q(n912) );
  hi1s1 U925 ( .DIN(n913), .Q(n600) );
  oai21s1 U926 ( .DIN1(n551), .DIN2(n914), .DIN3(n915), .Q(n913) );
  mxi21s1 U927 ( .DIN1(n916), .DIN2(n786), .SIN(N116), .Q(n915) );
  nor2s1 U928 ( .DIN1(N87), .DIN2(N107), .Q(n786) );
  nor2s1 U929 ( .DIN1(N87), .DIN2(n550), .Q(n916) );
  hi1s1 U930 ( .DIN(N107), .Q(n550) );
  xor2s1 U931 ( .DIN1(N116), .DIN2(N107), .Q(n914) );
  hi1s1 U932 ( .DIN(N87), .Q(n551) );
  xor2s1 U933 ( .DIN1(n917), .DIN2(n894), .Q(n782) );
  oai21s1 U934 ( .DIN1(n502), .DIN2(n513), .DIN3(n918), .Q(n894) );
  xor2s1 U935 ( .DIN1(n646), .DIN2(N77), .Q(n917) );
  hi1s1 U936 ( .DIN(N50), .Q(n646) );
  xnr2s1 U937 ( .DIN1(n678), .DIN2(n644), .Q(N323) );
  xnr2s1 U938 ( .DIN1(n919), .DIN2(n920), .Q(n644) );
  xnr2s1 U939 ( .DIN1(N244), .DIN2(n902), .Q(n920) );
  hi1s1 U940 ( .DIN(N238), .Q(n902) );
  xor2s1 U941 ( .DIN1(N226), .DIN2(n889), .Q(n919) );
  hi1s1 U942 ( .DIN(N232), .Q(n889) );
  xnr2s1 U943 ( .DIN1(n921), .DIN2(n922), .Q(n678) );
  xor2s1 U944 ( .DIN1(N257), .DIN2(N250), .Q(n922) );
  xnr2s1 U945 ( .DIN1(N270), .DIN2(N264), .Q(n921) );
  oai22s1 U946 ( .DIN1(n923), .DIN2(n924), .DIN3(n780), .DIN4(n925), .Q(N3195)
         );
  mxi21s1 U947 ( .DIN1(n781), .DIN2(n926), .SIN(n705), .Q(n925) );
  nnd2s1 U948 ( .DIN1(n783), .DIN2(N20), .Q(n705) );
  nor2s1 U949 ( .DIN1(n908), .DIN2(n683), .Q(n783) );
  hi1s1 U950 ( .DIN(N1), .Q(n683) );
  and4s1 U951 ( .DIN1(n927), .DIN2(n928), .DIN3(n929), .DIN4(n930), .Q(n926)
         );
  aoi22s1 U952 ( .DIN1(N264), .DIN2(N107), .DIN3(N270), .DIN4(N116), .Q(n930)
         );
  aoi22s1 U953 ( .DIN1(N226), .DIN2(N50), .DIN3(N232), .DIN4(N58), .Q(n929) );
  aoi22s1 U954 ( .DIN1(N238), .DIN2(N68), .DIN3(N244), .DIN4(N77), .Q(n928) );
  aoi22s1 U955 ( .DIN1(N250), .DIN2(N87), .DIN3(N257), .DIN4(N97), .Q(n927) );
  nnd2s1 U956 ( .DIN1(N50), .DIN2(n918), .Q(n781) );
  hi1s1 U957 ( .DIN(n780), .Q(n924) );
  nor2s1 U958 ( .DIN1(n682), .DIN2(n710), .Q(n780) );
  nnd2s1 U959 ( .DIN1(N1), .DIN2(n908), .Q(n710) );
  hi1s1 U960 ( .DIN(N13), .Q(n908) );
  hi1s1 U961 ( .DIN(N20), .Q(n682) );
  hi1s1 U962 ( .DIN(n931), .Q(n923) );
  oai21s1 U963 ( .DIN1(N257), .DIN2(N264), .DIN3(N250), .Q(n931) );
  nor3s1 U964 ( .DIN1(N50), .DIN2(N77), .DIN3(n918), .Q(N26) );
  nnd2s1 U965 ( .DIN1(n502), .DIN2(n513), .Q(n918) );
  hi1s1 U966 ( .DIN(N68), .Q(n513) );
  hi1s1 U967 ( .DIN(N58), .Q(n502) );
  oai21s1 U968 ( .DIN1(N97), .DIN2(N107), .DIN3(N87), .Q(N1947) );
endmodule

