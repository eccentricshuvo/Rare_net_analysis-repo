`timescale 1ns/10ps

module tb;
	reg N350;
	reg N349;
	reg N343;
	reg N330;
	reg N329;
	reg N326;
	reg N322;
	reg N317;
	reg N311;
	reg N303;
	reg N294;
	reg N283;
	reg N274;
	reg N270;
	reg N264;
	reg N257;
	reg N250;
	reg N244;
	reg N238;
	reg N232;
	reg N226;
	reg N223;
	reg N222;
	reg N213;
	reg N200;
	reg N190;
	reg N179;
	reg N169;
	reg N159;
	reg N150;
	reg N143;
	reg N137;
	reg N132;
	reg N128;
	reg N125;
	reg N124;
	reg N116;
	reg N107;
	reg N97;
	reg N87;
	reg N77;
	reg N68;
	reg N58;
	reg N50;
	reg N45;
	reg N41;
	reg N33;
	reg N20;
	reg N13;
	reg N1;
	wire N1713;
	wire N1947;
	wire N3195;
	wire N3833;
	wire N3987;
	wire N4028;
	wire N4145;
	wire N4589;
	wire N4667;
	wire N4815;
	wire N4944;
	wire N5002;
	wire N5045;
	wire N5047;
	wire N5078;
	wire N5102;
	wire N5120;
	wire N5121;
	wire N5192;
	wire N5231;
	wire N5360;
	wire N5361;

	c3540 uut(
		.N1(N1),
		.N13(N13),
		.N20(N20),
		.N33(N33),
		.N41(N41),
		.N45(N45),
		.N50(N50),
		.N58(N58),
		.N68(N68),
		.N77(N77),
		.N87(N87),
		.N97(N97),
		.N107(N107),
		.N116(N116),
		.N124(N124),
		.N125(N125),
		.N128(N128),
		.N132(N132),
		.N137(N137),
		.N143(N143),
		.N150(N150),
		.N159(N159),
		.N169(N169),
		.N179(N179),
		.N190(N190),
		.N200(N200),
		.N213(N213),
		.N222(N222),
		.N223(N223),
		.N226(N226),
		.N232(N232),
		.N238(N238),
		.N244(N244),
		.N250(N250),
		.N257(N257),
		.N264(N264),
		.N270(N270),
		.N274(N274),
		.N283(N283),
		.N294(N294),
		.N303(N303),
		.N311(N311),
		.N317(N317),
		.N322(N322),
		.N326(N326),
		.N329(N329),
		.N330(N330),
		.N343(N343),
		.N349(N349),
		.N350(N350),
		.N1713(N1713),
		.N1947(N1947),
		.N3195(N3195),
		.N3833(N3833),
		.N3987(N3987),
		.N4028(N4028),
		.N4145(N4145),
		.N4589(N4589),
		.N4667(N4667),
		.N4815(N4815),
		.N4944(N4944),
		.N5002(N5002),
		.N5045(N5045),
		.N5047(N5047),
		.N5078(N5078),
		.N5102(N5102),
		.N5120(N5120),
		.N5121(N5121),
		.N5192(N5192),
		.N5231(N5231),
		.N5360(N5360),
		.N5361(N5361)	);

	integer file, file_out;

	initial begin
		file_out=$fopen("./example/tb_log.txt");
		$dumpfile("output.vcd");
		$dumpvars(0,tb);
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = 0;
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = 50'b10011010100101101110010111110000101110100110110001;
		#10 $fwrite(file_out,"%b\n",{uut.N350,uut.N349,uut.N343,uut.N330,uut.N329,uut.N326,uut.N322,uut.N317,uut.N311,uut.N303,uut.N294,uut.N283,uut.N274,uut.N270,uut.N264,uut.N257,uut.N250,uut.N244,uut.N238,uut.N232,uut.N226,uut.N223,uut.N222,uut.N213,uut.N200,uut.N190,uut.N179,uut.N169,uut.N159,uut.N150,uut.N143,uut.N137,uut.N132,uut.N128,uut.N125,uut.N124,uut.N116,uut.N107,uut.N97,uut.N87,uut.N77,uut.N68,uut.N58,uut.N50,uut.N45,uut.N41,uut.N33,uut.N20,uut.N13,uut.N1,uut.N1713,uut.N1947,uut.N3195,uut.N3833,uut.N3987,uut.N4028,uut.N4145,uut.N4589,uut.N4667,uut.N4815,uut.N4944,uut.N5002,uut.N5045,uut.N5047,uut.N5078,uut.N5102,uut.N5120,uut.N5121,uut.N5192,uut.N5231,uut.N5360,uut.N5361,uut.n771,uut.N538,uut.n469,uut.n468,uut.n467,uut.n473,uut.n471,uut.n475,uut.n476,uut.n474,uut.n477,uut.n478,uut.n472,uut.n470,uut.n480,uut.n482,uut.n488,uut.n490,uut.n489,uut.n487,uut.n481,uut.n498,uut.n499,uut.n506,uut.n508,uut.n505,uut.n512,uut.n517,uut.n521,uut.n524,uut.n528,uut.n520,uut.n516,uut.n534,uut.n533,uut.n532,uut.n531,uut.N5080,uut.n540,uut.n542,uut.n541,uut.n545,uut.n549,uut.n548,uut.n547,uut.n546,uut.n544,uut.n557,uut.n560,uut.n561,uut.n556,uut.n555,uut.n539,uut.n567,uut.n507,uut.n511,uut.n566,uut.n570,uut.n543,uut.n574,uut.n581,uut.n584,uut.n585,uut.n587,uut.n591,uut.n590,uut.n589,uut.n588,uut.n586,uut.n595,uut.n594,uut.n593,uut.n592,uut.n583,uut.n582,uut.n599,uut.n578,uut.n602,uut.n603,uut.N5050,uut.n492,uut.n484,uut.n608,uut.n609,uut.n483,uut.n607,uut.n485,uut.n569,uut.n509,uut.n616,uut.n606,uut.n620,uut.n503,uut.n625,uut.n624,uut.n623,uut.n622,uut.n504,uut.n629,uut.n628,uut.n627,uut.n626,uut.n501,uut.n514,uut.n631,uut.n634,uut.n636,uut.n639,uut.n641,uut.n637,uut.n643,uut.n645,uut.n635,uut.n648,uut.n652,uut.n651,uut.n650,uut.n649,uut.n647,uut.n654,uut.n655,uut.n653,uut.n519,uut.n630,uut.n658,uut.n661,uut.n664,uut.n665,uut.n668,uut.n672,uut.n671,uut.n670,uut.n669,uut.n667,uut.n675,uut.n676,uut.n677,uut.n674,uut.n518,uut.n662,uut.n660,uut.n681,uut.n579,uut.n657,uut.n568,uut.n604,uut.n685,uut.n684,uut.n688,uut.n689,uut.n580,uut.n659,uut.n693,uut.n692,uut.n691,uut.n694,uut.n695,uut.n680,uut.n699,uut.n596,uut.n702,uut.n707,uut.n709,uut.n712,uut.n714,uut.n715,uut.n572,uut.n718,uut.n610,uut.n720,uut.n713,uut.n723,uut.n571,uut.n612,uut.n722,uut.n497,uut.n725,uut.n611,uut.n515,uut.n728,uut.n731,uut.n711,uut.n708,uut.n734,uut.n735,uut.n491,uut.n479,uut.n737,uut.n738,uut.n736,uut.n613,uut.n617,uut.n618,uut.n739,uut.n741,uut.n494,uut.n745,uut.n749,uut.n748,uut.n747,uut.n746,uut.n744,uut.n753,uut.n752,uut.n751,uut.n750,uut.n493,uut.n486,uut.n756,uut.n755,uut.n754,uut.n597,uut.n760,uut.n500,uut.n759,uut.n762,uut.n766,uut.n765,uut.n764,uut.n763,uut.n761,uut.n770,uut.n523,uut.n559,uut.n536,uut.n558,uut.n769,uut.n538,uut.n525,uut.n537,uut.n527,uut.n768,uut.n522,uut.n565,uut.n774,uut.n530,uut.n564,uut.n772,uut.n767,uut.n535,uut.n563,uut.n529,uut.n562,uut.n776,uut.n758,uut.n778,uut.n642,uut.n779,uut.n601,uut.n638,uut.n777,uut.n598,uut.n663,uut.n495,uut.n633,uut.n784,uut.n785,uut.n640,uut.n510,uut.n605,uut.n724,uut.n787,uut.n789,uut.n792,uut.n791,uut.n788,uut.n696,uut.n798,uut.n716,uut.n577,uut.n687,uut.n690,uut.n805,uut.n806,uut.n799,uut.n700,uut.n808,uut.n801,uut.n632,uut.n797,uut.n810,uut.n679,uut.n697,uut.n576,uut.n717,uut.n615,uut.n815,uut.n575,uut.n820,uut.n821,uut.n819,uut.n673,uut.n814,uut.n826,uut.n730,uut.n740,uut.n813,uut.n802,uut.n829,uut.n831,uut.n830,uut.n686,uut.n703,uut.n828,uut.n698,uut.n834,uut.n811,uut.n809,uut.n840,uut.n839,uut.n794,uut.n844,uut.n842,uut.n812,uut.n848,uut.n526,uut.n666,uut.n851,uut.n852,uut.n835,uut.n796,uut.n856,uut.n857,uut.n855,uut.n832,uut.n701,uut.n861,uut.n860,uut.n790,uut.n863,uut.n862,uut.n704,uut.n865,uut.n706,uut.n864,uut.n850,uut.n838,uut.n804,uut.n867,uut.n868,uut.n836,uut.n554,uut.n553,uut.n807,uut.n800,uut.n793,uut.n795,uut.n871,uut.n845,uut.n843,uut.n872,uut.n858,uut.n870,uut.n614,uut.n874,uut.n875,uut.n573,uut.n876,uut.n878,uut.n877,uut.n823,uut.n833,uut.n817,uut.n883,uut.n881,uut.n726,uut.n719,uut.n886,uut.n885,uut.n887,uut.n890,uut.n891,uut.n775,uut.n773,uut.n727,uut.n893,uut.n866,uut.n892,uut.n656,uut.n742,uut.n743,uut.n729,uut.n732,uut.n898,uut.n721,uut.n899,uut.n901,uut.n849,uut.n837,uut.n552,uut.n733,uut.n900,uut.n903,uut.n854,uut.n904,uut.n888,uut.n827,uut.n897,uut.n906,uut.n825,uut.n879,uut.n895,uut.n869,uut.n822,uut.n853,uut.n824,uut.n907,uut.n818,uut.n847,uut.n880,uut.n619,uut.n496,uut.n905,uut.n896,uut.n910,uut.n846,uut.n884,uut.n882,uut.n911,uut.n757,uut.n909,uut.n841,uut.n873,uut.n859,uut.n803,uut.n621,uut.n816,uut.n912,uut.n600,uut.n913,uut.n915,uut.n786,uut.n916,uut.n550,uut.n914,uut.n551,uut.n782,uut.n894,uut.n917,uut.n646,uut.N323,uut.n644,uut.n920,uut.n902,uut.n919,uut.n889,uut.n678,uut.n922,uut.n921,uut.n925,uut.n705,uut.n783,uut.n683,uut.n926,uut.n930,uut.n929,uut.n928,uut.n927,uut.n781,uut.n924,uut.n780,uut.n710,uut.n908,uut.n682,uut.n923,uut.n931,uut.N26,uut.n918,uut.n513,uut.n502});
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = 50'b10010010100101000000010011111110011011011101111110;
		#10 $fwrite(file_out,"%b\n",{uut.N350,uut.N349,uut.N343,uut.N330,uut.N329,uut.N326,uut.N322,uut.N317,uut.N311,uut.N303,uut.N294,uut.N283,uut.N274,uut.N270,uut.N264,uut.N257,uut.N250,uut.N244,uut.N238,uut.N232,uut.N226,uut.N223,uut.N222,uut.N213,uut.N200,uut.N190,uut.N179,uut.N169,uut.N159,uut.N150,uut.N143,uut.N137,uut.N132,uut.N128,uut.N125,uut.N124,uut.N116,uut.N107,uut.N97,uut.N87,uut.N77,uut.N68,uut.N58,uut.N50,uut.N45,uut.N41,uut.N33,uut.N20,uut.N13,uut.N1,uut.N1713,uut.N1947,uut.N3195,uut.N3833,uut.N3987,uut.N4028,uut.N4145,uut.N4589,uut.N4667,uut.N4815,uut.N4944,uut.N5002,uut.N5045,uut.N5047,uut.N5078,uut.N5102,uut.N5120,uut.N5121,uut.N5192,uut.N5231,uut.N5360,uut.N5361,uut.n771,uut.N538,uut.n469,uut.n468,uut.n467,uut.n473,uut.n471,uut.n475,uut.n476,uut.n474,uut.n477,uut.n478,uut.n472,uut.n470,uut.n480,uut.n482,uut.n488,uut.n490,uut.n489,uut.n487,uut.n481,uut.n498,uut.n499,uut.n506,uut.n508,uut.n505,uut.n512,uut.n517,uut.n521,uut.n524,uut.n528,uut.n520,uut.n516,uut.n534,uut.n533,uut.n532,uut.n531,uut.N5080,uut.n540,uut.n542,uut.n541,uut.n545,uut.n549,uut.n548,uut.n547,uut.n546,uut.n544,uut.n557,uut.n560,uut.n561,uut.n556,uut.n555,uut.n539,uut.n567,uut.n507,uut.n511,uut.n566,uut.n570,uut.n543,uut.n574,uut.n581,uut.n584,uut.n585,uut.n587,uut.n591,uut.n590,uut.n589,uut.n588,uut.n586,uut.n595,uut.n594,uut.n593,uut.n592,uut.n583,uut.n582,uut.n599,uut.n578,uut.n602,uut.n603,uut.N5050,uut.n492,uut.n484,uut.n608,uut.n609,uut.n483,uut.n607,uut.n485,uut.n569,uut.n509,uut.n616,uut.n606,uut.n620,uut.n503,uut.n625,uut.n624,uut.n623,uut.n622,uut.n504,uut.n629,uut.n628,uut.n627,uut.n626,uut.n501,uut.n514,uut.n631,uut.n634,uut.n636,uut.n639,uut.n641,uut.n637,uut.n643,uut.n645,uut.n635,uut.n648,uut.n652,uut.n651,uut.n650,uut.n649,uut.n647,uut.n654,uut.n655,uut.n653,uut.n519,uut.n630,uut.n658,uut.n661,uut.n664,uut.n665,uut.n668,uut.n672,uut.n671,uut.n670,uut.n669,uut.n667,uut.n675,uut.n676,uut.n677,uut.n674,uut.n518,uut.n662,uut.n660,uut.n681,uut.n579,uut.n657,uut.n568,uut.n604,uut.n685,uut.n684,uut.n688,uut.n689,uut.n580,uut.n659,uut.n693,uut.n692,uut.n691,uut.n694,uut.n695,uut.n680,uut.n699,uut.n596,uut.n702,uut.n707,uut.n709,uut.n712,uut.n714,uut.n715,uut.n572,uut.n718,uut.n610,uut.n720,uut.n713,uut.n723,uut.n571,uut.n612,uut.n722,uut.n497,uut.n725,uut.n611,uut.n515,uut.n728,uut.n731,uut.n711,uut.n708,uut.n734,uut.n735,uut.n491,uut.n479,uut.n737,uut.n738,uut.n736,uut.n613,uut.n617,uut.n618,uut.n739,uut.n741,uut.n494,uut.n745,uut.n749,uut.n748,uut.n747,uut.n746,uut.n744,uut.n753,uut.n752,uut.n751,uut.n750,uut.n493,uut.n486,uut.n756,uut.n755,uut.n754,uut.n597,uut.n760,uut.n500,uut.n759,uut.n762,uut.n766,uut.n765,uut.n764,uut.n763,uut.n761,uut.n770,uut.n523,uut.n559,uut.n536,uut.n558,uut.n769,uut.n538,uut.n525,uut.n537,uut.n527,uut.n768,uut.n522,uut.n565,uut.n774,uut.n530,uut.n564,uut.n772,uut.n767,uut.n535,uut.n563,uut.n529,uut.n562,uut.n776,uut.n758,uut.n778,uut.n642,uut.n779,uut.n601,uut.n638,uut.n777,uut.n598,uut.n663,uut.n495,uut.n633,uut.n784,uut.n785,uut.n640,uut.n510,uut.n605,uut.n724,uut.n787,uut.n789,uut.n792,uut.n791,uut.n788,uut.n696,uut.n798,uut.n716,uut.n577,uut.n687,uut.n690,uut.n805,uut.n806,uut.n799,uut.n700,uut.n808,uut.n801,uut.n632,uut.n797,uut.n810,uut.n679,uut.n697,uut.n576,uut.n717,uut.n615,uut.n815,uut.n575,uut.n820,uut.n821,uut.n819,uut.n673,uut.n814,uut.n826,uut.n730,uut.n740,uut.n813,uut.n802,uut.n829,uut.n831,uut.n830,uut.n686,uut.n703,uut.n828,uut.n698,uut.n834,uut.n811,uut.n809,uut.n840,uut.n839,uut.n794,uut.n844,uut.n842,uut.n812,uut.n848,uut.n526,uut.n666,uut.n851,uut.n852,uut.n835,uut.n796,uut.n856,uut.n857,uut.n855,uut.n832,uut.n701,uut.n861,uut.n860,uut.n790,uut.n863,uut.n862,uut.n704,uut.n865,uut.n706,uut.n864,uut.n850,uut.n838,uut.n804,uut.n867,uut.n868,uut.n836,uut.n554,uut.n553,uut.n807,uut.n800,uut.n793,uut.n795,uut.n871,uut.n845,uut.n843,uut.n872,uut.n858,uut.n870,uut.n614,uut.n874,uut.n875,uut.n573,uut.n876,uut.n878,uut.n877,uut.n823,uut.n833,uut.n817,uut.n883,uut.n881,uut.n726,uut.n719,uut.n886,uut.n885,uut.n887,uut.n890,uut.n891,uut.n775,uut.n773,uut.n727,uut.n893,uut.n866,uut.n892,uut.n656,uut.n742,uut.n743,uut.n729,uut.n732,uut.n898,uut.n721,uut.n899,uut.n901,uut.n849,uut.n837,uut.n552,uut.n733,uut.n900,uut.n903,uut.n854,uut.n904,uut.n888,uut.n827,uut.n897,uut.n906,uut.n825,uut.n879,uut.n895,uut.n869,uut.n822,uut.n853,uut.n824,uut.n907,uut.n818,uut.n847,uut.n880,uut.n619,uut.n496,uut.n905,uut.n896,uut.n910,uut.n846,uut.n884,uut.n882,uut.n911,uut.n757,uut.n909,uut.n841,uut.n873,uut.n859,uut.n803,uut.n621,uut.n816,uut.n912,uut.n600,uut.n913,uut.n915,uut.n786,uut.n916,uut.n550,uut.n914,uut.n551,uut.n782,uut.n894,uut.n917,uut.n646,uut.N323,uut.n644,uut.n920,uut.n902,uut.n919,uut.n889,uut.n678,uut.n922,uut.n921,uut.n925,uut.n705,uut.n783,uut.n683,uut.n926,uut.n930,uut.n929,uut.n928,uut.n927,uut.n781,uut.n924,uut.n780,uut.n710,uut.n908,uut.n682,uut.n923,uut.n931,uut.N26,uut.n918,uut.n513,uut.n502});
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = 50'b10010010100101101111000011100100110110001010110010;
		#10 $fwrite(file_out,"%b\n",{uut.N350,uut.N349,uut.N343,uut.N330,uut.N329,uut.N326,uut.N322,uut.N317,uut.N311,uut.N303,uut.N294,uut.N283,uut.N274,uut.N270,uut.N264,uut.N257,uut.N250,uut.N244,uut.N238,uut.N232,uut.N226,uut.N223,uut.N222,uut.N213,uut.N200,uut.N190,uut.N179,uut.N169,uut.N159,uut.N150,uut.N143,uut.N137,uut.N132,uut.N128,uut.N125,uut.N124,uut.N116,uut.N107,uut.N97,uut.N87,uut.N77,uut.N68,uut.N58,uut.N50,uut.N45,uut.N41,uut.N33,uut.N20,uut.N13,uut.N1,uut.N1713,uut.N1947,uut.N3195,uut.N3833,uut.N3987,uut.N4028,uut.N4145,uut.N4589,uut.N4667,uut.N4815,uut.N4944,uut.N5002,uut.N5045,uut.N5047,uut.N5078,uut.N5102,uut.N5120,uut.N5121,uut.N5192,uut.N5231,uut.N5360,uut.N5361,uut.n771,uut.N538,uut.n469,uut.n468,uut.n467,uut.n473,uut.n471,uut.n475,uut.n476,uut.n474,uut.n477,uut.n478,uut.n472,uut.n470,uut.n480,uut.n482,uut.n488,uut.n490,uut.n489,uut.n487,uut.n481,uut.n498,uut.n499,uut.n506,uut.n508,uut.n505,uut.n512,uut.n517,uut.n521,uut.n524,uut.n528,uut.n520,uut.n516,uut.n534,uut.n533,uut.n532,uut.n531,uut.N5080,uut.n540,uut.n542,uut.n541,uut.n545,uut.n549,uut.n548,uut.n547,uut.n546,uut.n544,uut.n557,uut.n560,uut.n561,uut.n556,uut.n555,uut.n539,uut.n567,uut.n507,uut.n511,uut.n566,uut.n570,uut.n543,uut.n574,uut.n581,uut.n584,uut.n585,uut.n587,uut.n591,uut.n590,uut.n589,uut.n588,uut.n586,uut.n595,uut.n594,uut.n593,uut.n592,uut.n583,uut.n582,uut.n599,uut.n578,uut.n602,uut.n603,uut.N5050,uut.n492,uut.n484,uut.n608,uut.n609,uut.n483,uut.n607,uut.n485,uut.n569,uut.n509,uut.n616,uut.n606,uut.n620,uut.n503,uut.n625,uut.n624,uut.n623,uut.n622,uut.n504,uut.n629,uut.n628,uut.n627,uut.n626,uut.n501,uut.n514,uut.n631,uut.n634,uut.n636,uut.n639,uut.n641,uut.n637,uut.n643,uut.n645,uut.n635,uut.n648,uut.n652,uut.n651,uut.n650,uut.n649,uut.n647,uut.n654,uut.n655,uut.n653,uut.n519,uut.n630,uut.n658,uut.n661,uut.n664,uut.n665,uut.n668,uut.n672,uut.n671,uut.n670,uut.n669,uut.n667,uut.n675,uut.n676,uut.n677,uut.n674,uut.n518,uut.n662,uut.n660,uut.n681,uut.n579,uut.n657,uut.n568,uut.n604,uut.n685,uut.n684,uut.n688,uut.n689,uut.n580,uut.n659,uut.n693,uut.n692,uut.n691,uut.n694,uut.n695,uut.n680,uut.n699,uut.n596,uut.n702,uut.n707,uut.n709,uut.n712,uut.n714,uut.n715,uut.n572,uut.n718,uut.n610,uut.n720,uut.n713,uut.n723,uut.n571,uut.n612,uut.n722,uut.n497,uut.n725,uut.n611,uut.n515,uut.n728,uut.n731,uut.n711,uut.n708,uut.n734,uut.n735,uut.n491,uut.n479,uut.n737,uut.n738,uut.n736,uut.n613,uut.n617,uut.n618,uut.n739,uut.n741,uut.n494,uut.n745,uut.n749,uut.n748,uut.n747,uut.n746,uut.n744,uut.n753,uut.n752,uut.n751,uut.n750,uut.n493,uut.n486,uut.n756,uut.n755,uut.n754,uut.n597,uut.n760,uut.n500,uut.n759,uut.n762,uut.n766,uut.n765,uut.n764,uut.n763,uut.n761,uut.n770,uut.n523,uut.n559,uut.n536,uut.n558,uut.n769,uut.n538,uut.n525,uut.n537,uut.n527,uut.n768,uut.n522,uut.n565,uut.n774,uut.n530,uut.n564,uut.n772,uut.n767,uut.n535,uut.n563,uut.n529,uut.n562,uut.n776,uut.n758,uut.n778,uut.n642,uut.n779,uut.n601,uut.n638,uut.n777,uut.n598,uut.n663,uut.n495,uut.n633,uut.n784,uut.n785,uut.n640,uut.n510,uut.n605,uut.n724,uut.n787,uut.n789,uut.n792,uut.n791,uut.n788,uut.n696,uut.n798,uut.n716,uut.n577,uut.n687,uut.n690,uut.n805,uut.n806,uut.n799,uut.n700,uut.n808,uut.n801,uut.n632,uut.n797,uut.n810,uut.n679,uut.n697,uut.n576,uut.n717,uut.n615,uut.n815,uut.n575,uut.n820,uut.n821,uut.n819,uut.n673,uut.n814,uut.n826,uut.n730,uut.n740,uut.n813,uut.n802,uut.n829,uut.n831,uut.n830,uut.n686,uut.n703,uut.n828,uut.n698,uut.n834,uut.n811,uut.n809,uut.n840,uut.n839,uut.n794,uut.n844,uut.n842,uut.n812,uut.n848,uut.n526,uut.n666,uut.n851,uut.n852,uut.n835,uut.n796,uut.n856,uut.n857,uut.n855,uut.n832,uut.n701,uut.n861,uut.n860,uut.n790,uut.n863,uut.n862,uut.n704,uut.n865,uut.n706,uut.n864,uut.n850,uut.n838,uut.n804,uut.n867,uut.n868,uut.n836,uut.n554,uut.n553,uut.n807,uut.n800,uut.n793,uut.n795,uut.n871,uut.n845,uut.n843,uut.n872,uut.n858,uut.n870,uut.n614,uut.n874,uut.n875,uut.n573,uut.n876,uut.n878,uut.n877,uut.n823,uut.n833,uut.n817,uut.n883,uut.n881,uut.n726,uut.n719,uut.n886,uut.n885,uut.n887,uut.n890,uut.n891,uut.n775,uut.n773,uut.n727,uut.n893,uut.n866,uut.n892,uut.n656,uut.n742,uut.n743,uut.n729,uut.n732,uut.n898,uut.n721,uut.n899,uut.n901,uut.n849,uut.n837,uut.n552,uut.n733,uut.n900,uut.n903,uut.n854,uut.n904,uut.n888,uut.n827,uut.n897,uut.n906,uut.n825,uut.n879,uut.n895,uut.n869,uut.n822,uut.n853,uut.n824,uut.n907,uut.n818,uut.n847,uut.n880,uut.n619,uut.n496,uut.n905,uut.n896,uut.n910,uut.n846,uut.n884,uut.n882,uut.n911,uut.n757,uut.n909,uut.n841,uut.n873,uut.n859,uut.n803,uut.n621,uut.n816,uut.n912,uut.n600,uut.n913,uut.n915,uut.n786,uut.n916,uut.n550,uut.n914,uut.n551,uut.n782,uut.n894,uut.n917,uut.n646,uut.N323,uut.n644,uut.n920,uut.n902,uut.n919,uut.n889,uut.n678,uut.n922,uut.n921,uut.n925,uut.n705,uut.n783,uut.n683,uut.n926,uut.n930,uut.n929,uut.n928,uut.n927,uut.n781,uut.n924,uut.n780,uut.n710,uut.n908,uut.n682,uut.n923,uut.n931,uut.N26,uut.n918,uut.n513,uut.n502});
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = 50'b10010010100101101111011100100001101010011000000100;
		#10 $fwrite(file_out,"%b\n",{uut.N350,uut.N349,uut.N343,uut.N330,uut.N329,uut.N326,uut.N322,uut.N317,uut.N311,uut.N303,uut.N294,uut.N283,uut.N274,uut.N270,uut.N264,uut.N257,uut.N250,uut.N244,uut.N238,uut.N232,uut.N226,uut.N223,uut.N222,uut.N213,uut.N200,uut.N190,uut.N179,uut.N169,uut.N159,uut.N150,uut.N143,uut.N137,uut.N132,uut.N128,uut.N125,uut.N124,uut.N116,uut.N107,uut.N97,uut.N87,uut.N77,uut.N68,uut.N58,uut.N50,uut.N45,uut.N41,uut.N33,uut.N20,uut.N13,uut.N1,uut.N1713,uut.N1947,uut.N3195,uut.N3833,uut.N3987,uut.N4028,uut.N4145,uut.N4589,uut.N4667,uut.N4815,uut.N4944,uut.N5002,uut.N5045,uut.N5047,uut.N5078,uut.N5102,uut.N5120,uut.N5121,uut.N5192,uut.N5231,uut.N5360,uut.N5361,uut.n771,uut.N538,uut.n469,uut.n468,uut.n467,uut.n473,uut.n471,uut.n475,uut.n476,uut.n474,uut.n477,uut.n478,uut.n472,uut.n470,uut.n480,uut.n482,uut.n488,uut.n490,uut.n489,uut.n487,uut.n481,uut.n498,uut.n499,uut.n506,uut.n508,uut.n505,uut.n512,uut.n517,uut.n521,uut.n524,uut.n528,uut.n520,uut.n516,uut.n534,uut.n533,uut.n532,uut.n531,uut.N5080,uut.n540,uut.n542,uut.n541,uut.n545,uut.n549,uut.n548,uut.n547,uut.n546,uut.n544,uut.n557,uut.n560,uut.n561,uut.n556,uut.n555,uut.n539,uut.n567,uut.n507,uut.n511,uut.n566,uut.n570,uut.n543,uut.n574,uut.n581,uut.n584,uut.n585,uut.n587,uut.n591,uut.n590,uut.n589,uut.n588,uut.n586,uut.n595,uut.n594,uut.n593,uut.n592,uut.n583,uut.n582,uut.n599,uut.n578,uut.n602,uut.n603,uut.N5050,uut.n492,uut.n484,uut.n608,uut.n609,uut.n483,uut.n607,uut.n485,uut.n569,uut.n509,uut.n616,uut.n606,uut.n620,uut.n503,uut.n625,uut.n624,uut.n623,uut.n622,uut.n504,uut.n629,uut.n628,uut.n627,uut.n626,uut.n501,uut.n514,uut.n631,uut.n634,uut.n636,uut.n639,uut.n641,uut.n637,uut.n643,uut.n645,uut.n635,uut.n648,uut.n652,uut.n651,uut.n650,uut.n649,uut.n647,uut.n654,uut.n655,uut.n653,uut.n519,uut.n630,uut.n658,uut.n661,uut.n664,uut.n665,uut.n668,uut.n672,uut.n671,uut.n670,uut.n669,uut.n667,uut.n675,uut.n676,uut.n677,uut.n674,uut.n518,uut.n662,uut.n660,uut.n681,uut.n579,uut.n657,uut.n568,uut.n604,uut.n685,uut.n684,uut.n688,uut.n689,uut.n580,uut.n659,uut.n693,uut.n692,uut.n691,uut.n694,uut.n695,uut.n680,uut.n699,uut.n596,uut.n702,uut.n707,uut.n709,uut.n712,uut.n714,uut.n715,uut.n572,uut.n718,uut.n610,uut.n720,uut.n713,uut.n723,uut.n571,uut.n612,uut.n722,uut.n497,uut.n725,uut.n611,uut.n515,uut.n728,uut.n731,uut.n711,uut.n708,uut.n734,uut.n735,uut.n491,uut.n479,uut.n737,uut.n738,uut.n736,uut.n613,uut.n617,uut.n618,uut.n739,uut.n741,uut.n494,uut.n745,uut.n749,uut.n748,uut.n747,uut.n746,uut.n744,uut.n753,uut.n752,uut.n751,uut.n750,uut.n493,uut.n486,uut.n756,uut.n755,uut.n754,uut.n597,uut.n760,uut.n500,uut.n759,uut.n762,uut.n766,uut.n765,uut.n764,uut.n763,uut.n761,uut.n770,uut.n523,uut.n559,uut.n536,uut.n558,uut.n769,uut.n538,uut.n525,uut.n537,uut.n527,uut.n768,uut.n522,uut.n565,uut.n774,uut.n530,uut.n564,uut.n772,uut.n767,uut.n535,uut.n563,uut.n529,uut.n562,uut.n776,uut.n758,uut.n778,uut.n642,uut.n779,uut.n601,uut.n638,uut.n777,uut.n598,uut.n663,uut.n495,uut.n633,uut.n784,uut.n785,uut.n640,uut.n510,uut.n605,uut.n724,uut.n787,uut.n789,uut.n792,uut.n791,uut.n788,uut.n696,uut.n798,uut.n716,uut.n577,uut.n687,uut.n690,uut.n805,uut.n806,uut.n799,uut.n700,uut.n808,uut.n801,uut.n632,uut.n797,uut.n810,uut.n679,uut.n697,uut.n576,uut.n717,uut.n615,uut.n815,uut.n575,uut.n820,uut.n821,uut.n819,uut.n673,uut.n814,uut.n826,uut.n730,uut.n740,uut.n813,uut.n802,uut.n829,uut.n831,uut.n830,uut.n686,uut.n703,uut.n828,uut.n698,uut.n834,uut.n811,uut.n809,uut.n840,uut.n839,uut.n794,uut.n844,uut.n842,uut.n812,uut.n848,uut.n526,uut.n666,uut.n851,uut.n852,uut.n835,uut.n796,uut.n856,uut.n857,uut.n855,uut.n832,uut.n701,uut.n861,uut.n860,uut.n790,uut.n863,uut.n862,uut.n704,uut.n865,uut.n706,uut.n864,uut.n850,uut.n838,uut.n804,uut.n867,uut.n868,uut.n836,uut.n554,uut.n553,uut.n807,uut.n800,uut.n793,uut.n795,uut.n871,uut.n845,uut.n843,uut.n872,uut.n858,uut.n870,uut.n614,uut.n874,uut.n875,uut.n573,uut.n876,uut.n878,uut.n877,uut.n823,uut.n833,uut.n817,uut.n883,uut.n881,uut.n726,uut.n719,uut.n886,uut.n885,uut.n887,uut.n890,uut.n891,uut.n775,uut.n773,uut.n727,uut.n893,uut.n866,uut.n892,uut.n656,uut.n742,uut.n743,uut.n729,uut.n732,uut.n898,uut.n721,uut.n899,uut.n901,uut.n849,uut.n837,uut.n552,uut.n733,uut.n900,uut.n903,uut.n854,uut.n904,uut.n888,uut.n827,uut.n897,uut.n906,uut.n825,uut.n879,uut.n895,uut.n869,uut.n822,uut.n853,uut.n824,uut.n907,uut.n818,uut.n847,uut.n880,uut.n619,uut.n496,uut.n905,uut.n896,uut.n910,uut.n846,uut.n884,uut.n882,uut.n911,uut.n757,uut.n909,uut.n841,uut.n873,uut.n859,uut.n803,uut.n621,uut.n816,uut.n912,uut.n600,uut.n913,uut.n915,uut.n786,uut.n916,uut.n550,uut.n914,uut.n551,uut.n782,uut.n894,uut.n917,uut.n646,uut.N323,uut.n644,uut.n920,uut.n902,uut.n919,uut.n889,uut.n678,uut.n922,uut.n921,uut.n925,uut.n705,uut.n783,uut.n683,uut.n926,uut.n930,uut.n929,uut.n928,uut.n927,uut.n781,uut.n924,uut.n780,uut.n710,uut.n908,uut.n682,uut.n923,uut.n931,uut.N26,uut.n918,uut.n513,uut.n502});
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = 50'b10011010100101100000111111100000011110110000001100;
		#10 $fwrite(file_out,"%b\n",{uut.N350,uut.N349,uut.N343,uut.N330,uut.N329,uut.N326,uut.N322,uut.N317,uut.N311,uut.N303,uut.N294,uut.N283,uut.N274,uut.N270,uut.N264,uut.N257,uut.N250,uut.N244,uut.N238,uut.N232,uut.N226,uut.N223,uut.N222,uut.N213,uut.N200,uut.N190,uut.N179,uut.N169,uut.N159,uut.N150,uut.N143,uut.N137,uut.N132,uut.N128,uut.N125,uut.N124,uut.N116,uut.N107,uut.N97,uut.N87,uut.N77,uut.N68,uut.N58,uut.N50,uut.N45,uut.N41,uut.N33,uut.N20,uut.N13,uut.N1,uut.N1713,uut.N1947,uut.N3195,uut.N3833,uut.N3987,uut.N4028,uut.N4145,uut.N4589,uut.N4667,uut.N4815,uut.N4944,uut.N5002,uut.N5045,uut.N5047,uut.N5078,uut.N5102,uut.N5120,uut.N5121,uut.N5192,uut.N5231,uut.N5360,uut.N5361,uut.n771,uut.N538,uut.n469,uut.n468,uut.n467,uut.n473,uut.n471,uut.n475,uut.n476,uut.n474,uut.n477,uut.n478,uut.n472,uut.n470,uut.n480,uut.n482,uut.n488,uut.n490,uut.n489,uut.n487,uut.n481,uut.n498,uut.n499,uut.n506,uut.n508,uut.n505,uut.n512,uut.n517,uut.n521,uut.n524,uut.n528,uut.n520,uut.n516,uut.n534,uut.n533,uut.n532,uut.n531,uut.N5080,uut.n540,uut.n542,uut.n541,uut.n545,uut.n549,uut.n548,uut.n547,uut.n546,uut.n544,uut.n557,uut.n560,uut.n561,uut.n556,uut.n555,uut.n539,uut.n567,uut.n507,uut.n511,uut.n566,uut.n570,uut.n543,uut.n574,uut.n581,uut.n584,uut.n585,uut.n587,uut.n591,uut.n590,uut.n589,uut.n588,uut.n586,uut.n595,uut.n594,uut.n593,uut.n592,uut.n583,uut.n582,uut.n599,uut.n578,uut.n602,uut.n603,uut.N5050,uut.n492,uut.n484,uut.n608,uut.n609,uut.n483,uut.n607,uut.n485,uut.n569,uut.n509,uut.n616,uut.n606,uut.n620,uut.n503,uut.n625,uut.n624,uut.n623,uut.n622,uut.n504,uut.n629,uut.n628,uut.n627,uut.n626,uut.n501,uut.n514,uut.n631,uut.n634,uut.n636,uut.n639,uut.n641,uut.n637,uut.n643,uut.n645,uut.n635,uut.n648,uut.n652,uut.n651,uut.n650,uut.n649,uut.n647,uut.n654,uut.n655,uut.n653,uut.n519,uut.n630,uut.n658,uut.n661,uut.n664,uut.n665,uut.n668,uut.n672,uut.n671,uut.n670,uut.n669,uut.n667,uut.n675,uut.n676,uut.n677,uut.n674,uut.n518,uut.n662,uut.n660,uut.n681,uut.n579,uut.n657,uut.n568,uut.n604,uut.n685,uut.n684,uut.n688,uut.n689,uut.n580,uut.n659,uut.n693,uut.n692,uut.n691,uut.n694,uut.n695,uut.n680,uut.n699,uut.n596,uut.n702,uut.n707,uut.n709,uut.n712,uut.n714,uut.n715,uut.n572,uut.n718,uut.n610,uut.n720,uut.n713,uut.n723,uut.n571,uut.n612,uut.n722,uut.n497,uut.n725,uut.n611,uut.n515,uut.n728,uut.n731,uut.n711,uut.n708,uut.n734,uut.n735,uut.n491,uut.n479,uut.n737,uut.n738,uut.n736,uut.n613,uut.n617,uut.n618,uut.n739,uut.n741,uut.n494,uut.n745,uut.n749,uut.n748,uut.n747,uut.n746,uut.n744,uut.n753,uut.n752,uut.n751,uut.n750,uut.n493,uut.n486,uut.n756,uut.n755,uut.n754,uut.n597,uut.n760,uut.n500,uut.n759,uut.n762,uut.n766,uut.n765,uut.n764,uut.n763,uut.n761,uut.n770,uut.n523,uut.n559,uut.n536,uut.n558,uut.n769,uut.n538,uut.n525,uut.n537,uut.n527,uut.n768,uut.n522,uut.n565,uut.n774,uut.n530,uut.n564,uut.n772,uut.n767,uut.n535,uut.n563,uut.n529,uut.n562,uut.n776,uut.n758,uut.n778,uut.n642,uut.n779,uut.n601,uut.n638,uut.n777,uut.n598,uut.n663,uut.n495,uut.n633,uut.n784,uut.n785,uut.n640,uut.n510,uut.n605,uut.n724,uut.n787,uut.n789,uut.n792,uut.n791,uut.n788,uut.n696,uut.n798,uut.n716,uut.n577,uut.n687,uut.n690,uut.n805,uut.n806,uut.n799,uut.n700,uut.n808,uut.n801,uut.n632,uut.n797,uut.n810,uut.n679,uut.n697,uut.n576,uut.n717,uut.n615,uut.n815,uut.n575,uut.n820,uut.n821,uut.n819,uut.n673,uut.n814,uut.n826,uut.n730,uut.n740,uut.n813,uut.n802,uut.n829,uut.n831,uut.n830,uut.n686,uut.n703,uut.n828,uut.n698,uut.n834,uut.n811,uut.n809,uut.n840,uut.n839,uut.n794,uut.n844,uut.n842,uut.n812,uut.n848,uut.n526,uut.n666,uut.n851,uut.n852,uut.n835,uut.n796,uut.n856,uut.n857,uut.n855,uut.n832,uut.n701,uut.n861,uut.n860,uut.n790,uut.n863,uut.n862,uut.n704,uut.n865,uut.n706,uut.n864,uut.n850,uut.n838,uut.n804,uut.n867,uut.n868,uut.n836,uut.n554,uut.n553,uut.n807,uut.n800,uut.n793,uut.n795,uut.n871,uut.n845,uut.n843,uut.n872,uut.n858,uut.n870,uut.n614,uut.n874,uut.n875,uut.n573,uut.n876,uut.n878,uut.n877,uut.n823,uut.n833,uut.n817,uut.n883,uut.n881,uut.n726,uut.n719,uut.n886,uut.n885,uut.n887,uut.n890,uut.n891,uut.n775,uut.n773,uut.n727,uut.n893,uut.n866,uut.n892,uut.n656,uut.n742,uut.n743,uut.n729,uut.n732,uut.n898,uut.n721,uut.n899,uut.n901,uut.n849,uut.n837,uut.n552,uut.n733,uut.n900,uut.n903,uut.n854,uut.n904,uut.n888,uut.n827,uut.n897,uut.n906,uut.n825,uut.n879,uut.n895,uut.n869,uut.n822,uut.n853,uut.n824,uut.n907,uut.n818,uut.n847,uut.n880,uut.n619,uut.n496,uut.n905,uut.n896,uut.n910,uut.n846,uut.n884,uut.n882,uut.n911,uut.n757,uut.n909,uut.n841,uut.n873,uut.n859,uut.n803,uut.n621,uut.n816,uut.n912,uut.n600,uut.n913,uut.n915,uut.n786,uut.n916,uut.n550,uut.n914,uut.n551,uut.n782,uut.n894,uut.n917,uut.n646,uut.N323,uut.n644,uut.n920,uut.n902,uut.n919,uut.n889,uut.n678,uut.n922,uut.n921,uut.n925,uut.n705,uut.n783,uut.n683,uut.n926,uut.n930,uut.n929,uut.n928,uut.n927,uut.n781,uut.n924,uut.n780,uut.n710,uut.n908,uut.n682,uut.n923,uut.n931,uut.N26,uut.n918,uut.n513,uut.n502});
		{N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350} = 50'b10011010100101100010000011000000011111010100101100;
		#10 $fwrite(file_out,"%b\n",{uut.N350,uut.N349,uut.N343,uut.N330,uut.N329,uut.N326,uut.N322,uut.N317,uut.N311,uut.N303,uut.N294,uut.N283,uut.N274,uut.N270,uut.N264,uut.N257,uut.N250,uut.N244,uut.N238,uut.N232,uut.N226,uut.N223,uut.N222,uut.N213,uut.N200,uut.N190,uut.N179,uut.N169,uut.N159,uut.N150,uut.N143,uut.N137,uut.N132,uut.N128,uut.N125,uut.N124,uut.N116,uut.N107,uut.N97,uut.N87,uut.N77,uut.N68,uut.N58,uut.N50,uut.N45,uut.N41,uut.N33,uut.N20,uut.N13,uut.N1,uut.N1713,uut.N1947,uut.N3195,uut.N3833,uut.N3987,uut.N4028,uut.N4145,uut.N4589,uut.N4667,uut.N4815,uut.N4944,uut.N5002,uut.N5045,uut.N5047,uut.N5078,uut.N5102,uut.N5120,uut.N5121,uut.N5192,uut.N5231,uut.N5360,uut.N5361,uut.n771,uut.N538,uut.n469,uut.n468,uut.n467,uut.n473,uut.n471,uut.n475,uut.n476,uut.n474,uut.n477,uut.n478,uut.n472,uut.n470,uut.n480,uut.n482,uut.n488,uut.n490,uut.n489,uut.n487,uut.n481,uut.n498,uut.n499,uut.n506,uut.n508,uut.n505,uut.n512,uut.n517,uut.n521,uut.n524,uut.n528,uut.n520,uut.n516,uut.n534,uut.n533,uut.n532,uut.n531,uut.N5080,uut.n540,uut.n542,uut.n541,uut.n545,uut.n549,uut.n548,uut.n547,uut.n546,uut.n544,uut.n557,uut.n560,uut.n561,uut.n556,uut.n555,uut.n539,uut.n567,uut.n507,uut.n511,uut.n566,uut.n570,uut.n543,uut.n574,uut.n581,uut.n584,uut.n585,uut.n587,uut.n591,uut.n590,uut.n589,uut.n588,uut.n586,uut.n595,uut.n594,uut.n593,uut.n592,uut.n583,uut.n582,uut.n599,uut.n578,uut.n602,uut.n603,uut.N5050,uut.n492,uut.n484,uut.n608,uut.n609,uut.n483,uut.n607,uut.n485,uut.n569,uut.n509,uut.n616,uut.n606,uut.n620,uut.n503,uut.n625,uut.n624,uut.n623,uut.n622,uut.n504,uut.n629,uut.n628,uut.n627,uut.n626,uut.n501,uut.n514,uut.n631,uut.n634,uut.n636,uut.n639,uut.n641,uut.n637,uut.n643,uut.n645,uut.n635,uut.n648,uut.n652,uut.n651,uut.n650,uut.n649,uut.n647,uut.n654,uut.n655,uut.n653,uut.n519,uut.n630,uut.n658,uut.n661,uut.n664,uut.n665,uut.n668,uut.n672,uut.n671,uut.n670,uut.n669,uut.n667,uut.n675,uut.n676,uut.n677,uut.n674,uut.n518,uut.n662,uut.n660,uut.n681,uut.n579,uut.n657,uut.n568,uut.n604,uut.n685,uut.n684,uut.n688,uut.n689,uut.n580,uut.n659,uut.n693,uut.n692,uut.n691,uut.n694,uut.n695,uut.n680,uut.n699,uut.n596,uut.n702,uut.n707,uut.n709,uut.n712,uut.n714,uut.n715,uut.n572,uut.n718,uut.n610,uut.n720,uut.n713,uut.n723,uut.n571,uut.n612,uut.n722,uut.n497,uut.n725,uut.n611,uut.n515,uut.n728,uut.n731,uut.n711,uut.n708,uut.n734,uut.n735,uut.n491,uut.n479,uut.n737,uut.n738,uut.n736,uut.n613,uut.n617,uut.n618,uut.n739,uut.n741,uut.n494,uut.n745,uut.n749,uut.n748,uut.n747,uut.n746,uut.n744,uut.n753,uut.n752,uut.n751,uut.n750,uut.n493,uut.n486,uut.n756,uut.n755,uut.n754,uut.n597,uut.n760,uut.n500,uut.n759,uut.n762,uut.n766,uut.n765,uut.n764,uut.n763,uut.n761,uut.n770,uut.n523,uut.n559,uut.n536,uut.n558,uut.n769,uut.n538,uut.n525,uut.n537,uut.n527,uut.n768,uut.n522,uut.n565,uut.n774,uut.n530,uut.n564,uut.n772,uut.n767,uut.n535,uut.n563,uut.n529,uut.n562,uut.n776,uut.n758,uut.n778,uut.n642,uut.n779,uut.n601,uut.n638,uut.n777,uut.n598,uut.n663,uut.n495,uut.n633,uut.n784,uut.n785,uut.n640,uut.n510,uut.n605,uut.n724,uut.n787,uut.n789,uut.n792,uut.n791,uut.n788,uut.n696,uut.n798,uut.n716,uut.n577,uut.n687,uut.n690,uut.n805,uut.n806,uut.n799,uut.n700,uut.n808,uut.n801,uut.n632,uut.n797,uut.n810,uut.n679,uut.n697,uut.n576,uut.n717,uut.n615,uut.n815,uut.n575,uut.n820,uut.n821,uut.n819,uut.n673,uut.n814,uut.n826,uut.n730,uut.n740,uut.n813,uut.n802,uut.n829,uut.n831,uut.n830,uut.n686,uut.n703,uut.n828,uut.n698,uut.n834,uut.n811,uut.n809,uut.n840,uut.n839,uut.n794,uut.n844,uut.n842,uut.n812,uut.n848,uut.n526,uut.n666,uut.n851,uut.n852,uut.n835,uut.n796,uut.n856,uut.n857,uut.n855,uut.n832,uut.n701,uut.n861,uut.n860,uut.n790,uut.n863,uut.n862,uut.n704,uut.n865,uut.n706,uut.n864,uut.n850,uut.n838,uut.n804,uut.n867,uut.n868,uut.n836,uut.n554,uut.n553,uut.n807,uut.n800,uut.n793,uut.n795,uut.n871,uut.n845,uut.n843,uut.n872,uut.n858,uut.n870,uut.n614,uut.n874,uut.n875,uut.n573,uut.n876,uut.n878,uut.n877,uut.n823,uut.n833,uut.n817,uut.n883,uut.n881,uut.n726,uut.n719,uut.n886,uut.n885,uut.n887,uut.n890,uut.n891,uut.n775,uut.n773,uut.n727,uut.n893,uut.n866,uut.n892,uut.n656,uut.n742,uut.n743,uut.n729,uut.n732,uut.n898,uut.n721,uut.n899,uut.n901,uut.n849,uut.n837,uut.n552,uut.n733,uut.n900,uut.n903,uut.n854,uut.n904,uut.n888,uut.n827,uut.n897,uut.n906,uut.n825,uut.n879,uut.n895,uut.n869,uut.n822,uut.n853,uut.n824,uut.n907,uut.n818,uut.n847,uut.n880,uut.n619,uut.n496,uut.n905,uut.n896,uut.n910,uut.n846,uut.n884,uut.n882,uut.n911,uut.n757,uut.n909,uut.n841,uut.n873,uut.n859,uut.n803,uut.n621,uut.n816,uut.n912,uut.n600,uut.n913,uut.n915,uut.n786,uut.n916,uut.n550,uut.n914,uut.n551,uut.n782,uut.n894,uut.n917,uut.n646,uut.N323,uut.n644,uut.n920,uut.n902,uut.n919,uut.n889,uut.n678,uut.n922,uut.n921,uut.n925,uut.n705,uut.n783,uut.n683,uut.n926,uut.n930,uut.n929,uut.n928,uut.n927,uut.n781,uut.n924,uut.n780,uut.n710,uut.n908,uut.n682,uut.n923,uut.n931,uut.N26,uut.n918,uut.n513,uut.n502});
		#100 $finish;
	end
endmodule